* Copyright 2025 ICsprout Integrated Circuit Co., Ltd.
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

************************************************************************
* Library Name: ICSCORE
* Cell Name:    INV
* View Name:    schematic
************************************************************************

.SUBCKT INV A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MMN0 Y A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    ADDFX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT ADDFX1H7L A B CI CO S VDD VSS
*.PININFO A:I B:I CI:I CO:O S:O VDD:B VSS:B
MMM12 net90 A net29 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM10 net29 net62 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM2 net9 B VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM11 net90 B net29 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM6 net25 CI VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM13 net90 CI net29 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM7 net62 A net25 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM8 net62 B net25 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM25 net49 B VDD VDD pm1p2_lvt_lp W=230n L=60n m=1
MMM23 net90 A net53 VDD pm1p2_lvt_lp W=230n L=60n m=1
MMM0 net62 A net9 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM22 net53 CI net49 VDD pm1p2_lvt_lp W=230n L=60n m=1
MMM20 net102 CI net110 VSS nm1p2_lvt_lp W=180n L=60n m=1
MMM3 net66 B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM24 net110 B VSS VSS nm1p2_lvt_lp W=180n L=60n m=1
MMM5 net62 A net77 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM14 net93 net62 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM16 net90 A net93 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM1 net62 A net66 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM17 net90 CI net93 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM15 net90 B net93 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM9 net62 B net77 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM21 net90 A net102 VSS nm1p2_lvt_lp W=180n L=60n m=1
MMM4 net77 CI VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
XI2 net90 VDD VSS S / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
XXI2 net62 VDD VSS CO / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    ADDFX1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT ADDFX1P4H7L A B CI CO S VDD VSS
*.PININFO A:I B:I CI:I CO:O S:O VDD:B VSS:B
MMM12 net90 A net29 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM10 net29 net62 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM2 net9 B VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM11 net90 B net29 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM6 net25 CI VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM13 net90 CI net29 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM7 net62 A net25 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM8 net62 B net25 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM25 net49 B VDD VDD pm1p2_lvt_lp W=230n L=60n m=1
MMM23 net90 A net53 VDD pm1p2_lvt_lp W=230n L=60n m=1
MMM0 net62 A net9 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM22 net53 CI net49 VDD pm1p2_lvt_lp W=230n L=60n m=1
MMM20 net102 CI net110 VSS nm1p2_lvt_lp W=180n L=60n m=1
MMM3 net66 B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM24 net110 B VSS VSS nm1p2_lvt_lp W=180n L=60n m=1
MMM5 net62 A net77 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM14 net93 net62 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM16 net90 A net93 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM1 net62 A net66 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM17 net90 CI net93 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM15 net90 B net93 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM9 net62 B net77 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM21 net90 A net102 VSS nm1p2_lvt_lp W=180n L=60n m=1
MMM4 net77 CI VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
XI3 net90 VDD VSS S / INV pl=6e-08 pw=3.14e-07 nl=6e-08 nw=2.46e-07
XXI2 net62 VDD VSS CO / INV pl=6e-08 pw=3.14e-07 nl=6e-08 nw=2.46e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    ADDFX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT ADDFX2H7L A B CI CO S VDD VSS
*.PININFO A:I B:I CI:I CO:O S:O VDD:B VSS:B
XI14 net30 VDD VSS S / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
XXI2 net58 VDD VSS CO / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
MMM17 net30 CI net33 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM16 net30 A net33 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM24 net10 B VSS VSS nm1p2_lvt_lp W=180n L=60n m=1
MMM15 net30 B net33 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM20 net18 CI net10 VSS nm1p2_lvt_lp W=180n L=60n m=1
MMM14 net33 net58 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM9 net58 B net49 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM21 net30 A net18 VSS nm1p2_lvt_lp W=180n L=60n m=1
MMM5 net58 A net49 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM1 net58 A net54 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM3 net54 B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM4 net49 CI VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM6 net101 CI VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM25 net77 B VDD VDD pm1p2_lvt_lp W=230n L=60n m=1
MMM2 net117 B VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM22 net73 CI net77 VDD pm1p2_lvt_lp W=230n L=60n m=1
MMM13 net30 CI net97 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM10 net97 net58 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM7 net58 A net101 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM12 net30 A net97 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM11 net30 B net97 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM0 net58 A net117 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM8 net58 B net101 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM23 net30 A net73 VDD pm1p2_lvt_lp W=230n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net15 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 net15 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP2 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    ADDHX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT ADDHX1H7L A B CO S VDD VSS
*.PININFO A:I B:I CO:O S:O VDD:B VSS:B
XI13 BN B net45 net_25 VDD VSS / TG pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI12 B BN net034 net_25 VDD VSS / TG pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI12 A VDD VSS net45 / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI14 net_25 VDD VSS S / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI11 net45 VDD VSS net034 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI9 B VDD VSS BN / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI11 net_7 VDD VSS CO / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI10 B A VDD VSS net_7 / NAND2 pl=6E-08 pw=2E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net15 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 net15 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP2 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    ADDHX1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT ADDHX1P4H7L A B CO S VDD VSS
*.PININFO A:I B:I CO:O S:O VDD:B VSS:B
XI18 BN B net45 net_25 VDD VSS / TG pl=6E-08 pw=3.64E-07 nl=6E-08 nw=2.56E-07
XI9 B BN net034 net_25 VDD VSS / TG pl=6E-08 pw=3.64E-07 nl=6E-08 nw=2.56E-07
XI20 A VDD VSS net45 / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI15 net_25 VDD VSS S / INV pl=6E-08 pw=3.64E-07 nl=6E-08 nw=2.56E-07
XI17 B VDD VSS BN / INV pl=6E-08 pw=3.64E-07 nl=6E-08 nw=2.56E-07
XI16 net45 VDD VSS net034 / INV pl=6E-08 pw=3.64E-07 nl=6E-08 nw=2.56E-07
XI19 net_7 VDD VSS CO / INV pl=6E-08 pw=3.64E-07 nl=6E-08 nw=2.56E-07
XI11 B A VDD VSS net_7 / NAND2 pl=6E-08 pw=2E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net15 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 net15 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP2 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    ADDHX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT ADDHX2H7L A B CO S VDD VSS
*.PININFO A:I B:I CO:O S:O VDD:B VSS:B
XI14 BN B net45 net_25 VDD VSS / TG pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI9 B BN net034 net_25 VDD VSS / TG pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI8 A VDD VSS net45 / INV pl=6E-08 pw=6E-07 nl=6E-08 nw=4.2E-07
XI15 net_25 VDD VSS S / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI13 net45 VDD VSS net034 / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI10 B VDD VSS BN / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI12 net_7 VDD VSS CO / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI11 B A VDD VSS net_7 / NAND2 pl=6E-08 pw=2E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND2X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND2X0P5H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 net26 B net6 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 net6 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP1 net26 B VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP0 net26 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI2 net26 VDD VSS Y / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND2X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND2X0P7H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 net26 B net6 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 net6 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP1 net26 B VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP0 net26 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI2 net26 VDD VSS Y / INV pl=6e-08 pw=2.22e-07 nl=6e-08 nw=1.74e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND2X12H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND2X12H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 net26 B net6 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN1 net6 A VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMP1 net26 B VDD VDD pm1p2_lvt_lp W=930n L=60n m=1
MMP0 net26 A VDD VDD pm1p2_lvt_lp W=930n L=60n m=1
XXI2 net26 VDD VSS Y / INV pl=6e-08 pw=22.8e-07 nl=6e-08 nw=18e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND2X16H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND2X16H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 net26 B net6 VSS nm1p2_lvt_lp W=1.2u L=60n m=1
MMN1 net6 A VSS VSS nm1p2_lvt_lp W=1.2u L=60n m=1
MMP1 net26 B VDD VDD pm1p2_lvt_lp W=1.24u L=60n m=1
MMP0 net26 A VDD VDD pm1p2_lvt_lp W=1.24u L=60n m=1
XXI2 net26 VDD VSS Y / INV pl=6e-08 pw=30.4e-07 nl=6e-08 nw=24e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND2X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND2X1H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 net26 B net6 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 net6 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM0 net26 B VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP0 net26 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI2 net26 VDD VSS Y / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND2X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND2X1P4H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 net26 B net6 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 net6 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP1 net26 B VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP0 net26 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI2 net26 VDD VSS Y / INV pl=6e-08 pw=3.14e-07 nl=6e-08 nw=2.46e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND2X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND2X2H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 net26 B net6 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 net6 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP1 net26 B VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP0 net26 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI2 net26 VDD VSS Y / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND2X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND2X3H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 net26 B net6 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 net6 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP1 net26 B VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP0 net26 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI2 net26 VDD VSS Y / INV pl=6e-08 pw=5.7e-07 nl=6e-08 nw=4.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND2X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND2X4H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 net26 B net6 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN1 net6 A VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP1 net26 B VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MMP0 net26 A VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
XXI2 net26 VDD VSS Y / INV pl=6e-08 pw=7.6e-07 nl=6e-08 nw=6e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND2X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND2X6H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 net26 B net6 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN1 net6 A VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP1 net26 B VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP0 net26 A VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
XXI2 net26 VDD VSS Y / INV pl=6e-08 pw=11.4e-07 nl=6e-08 nw=9e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND2X8H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND2X8H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 net26 B net6 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN1 net6 A VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMP1 net26 B VDD VDD pm1p2_lvt_lp W=620n L=60n m=1
MMP0 net26 A VDD VDD pm1p2_lvt_lp W=620n L=60n m=1
XXI2 net26 VDD VSS Y / INV pl=6e-08 pw=15.2e-07 nl=6e-08 nw=12e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND3X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND3X0P5H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN0 net36 C net10 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net7 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP0 net36 A VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net36 B VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP2 net36 C VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
XI0 net36 VDD VSS Y / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND3X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND3X0P7H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net7 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 net36 C net10 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP2 net36 C VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net36 B VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP0 net36 A VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
XI1 net36 VDD VSS Y / INV pl=6e-08 pw=2.22e-07 nl=6e-08 nw=1.74e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND3X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND3X1H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net7 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 net36 C net10 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP2 net36 C VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net36 B VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP0 net36 A VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
XI1 net36 VDD VSS Y / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND3X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND3X1P4H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net7 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 net36 C net10 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP2 net36 C VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net36 B VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP0 net36 A VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
XI1 net36 VDD VSS Y / INV pl=6e-08 pw=3.14e-07 nl=6e-08 nw=2.46e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND3X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND3X2H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN0 net36 C net10 VSS nm1p2_lvt_lp W=160n L=60n m=1
MMN4 net7 A VSS VSS nm1p2_lvt_lp W=160n L=60n m=1
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=160n L=60n m=1
MMP0 net36 A VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net36 B VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP2 net36 C VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
XI0 net36 VDD VSS Y / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND3X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND3X3H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net7 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 net36 C net10 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP2 net36 C VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 net36 B VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP0 net36 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XI1 net36 VDD VSS Y / INV pl=6e-08 pw=5.7e-07 nl=6e-08 nw=4.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND3X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND3X4H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN0 net36 C net10 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN4 net7 A VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP0 net36 A VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP1 net36 B VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP2 net36 C VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
XI0 net36 VDD VSS Y / INV pl=6e-08 pw=7.6e-07 nl=6e-08 nw=6e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND3X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND3X6H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN0 net36 C net10 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN4 net7 A VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP0 net36 A VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP1 net36 B VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP2 net36 C VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
XI0 net36 VDD VSS Y / INV pl=6e-08 pw=11.4e-07 nl=6e-08 nw=9e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND3X8H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND3X8H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN0 net36 C net10 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN4 net7 A VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMP0 net36 A VDD VDD pm1p2_lvt_lp W=540n L=60n m=1
MMP1 net36 B VDD VDD pm1p2_lvt_lp W=540n L=60n m=1
MMP2 net36 C VDD VDD pm1p2_lvt_lp W=540n L=60n m=1
XI0 net36 VDD VSS Y / INV pl=6e-08 pw=15.2e-07 nl=6e-08 nw=12e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND4X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND4X0P5H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MNM0 net35 D net45 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net45 C net42 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 net42 B net39 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM3 net39 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM0 net35 A VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM1 net35 B VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM2 net35 C VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM3 net35 D VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
XI0 net35 VDD VSS Y / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND4X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND4X0P7H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MNM0 net35 D net45 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net45 C net42 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 net42 B net39 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM3 net39 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM0 net35 A VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM1 net35 B VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM2 net35 C VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM3 net35 D VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
XI0 net35 VDD VSS Y / INV pl=6e-08 pw=2.22e-07 nl=6e-08 nw=1.74e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND4X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND4X1H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 B net28 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net28 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 net35 D net10 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP3 net35 A VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP2 net35 D VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net35 C VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP0 net35 B VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
XXI2 net35 VDD VSS Y / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND4X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND4X1P4H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MNM0 net35 D net45 VSS nm1p2_lvt_lp W=160n L=60n m=1
MNM1 net45 C net42 VSS nm1p2_lvt_lp W=160n L=60n m=1
MNM2 net42 B net39 VSS nm1p2_lvt_lp W=160n L=60n m=1
MNM3 net39 A VSS VSS nm1p2_lvt_lp W=160n L=60n m=1
MPM0 net35 A VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM1 net35 B VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM2 net35 C VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM3 net35 D VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
XI0 net35 VDD VSS Y / INV pl=6e-08 pw=3.14e-07 nl=6e-08 nw=2.46e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND4X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND4X2H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MNM4 net35 D net45 VSS nm1p2_lvt_lp W=170n L=60n m=1
MNM5 net45 C net42 VSS nm1p2_lvt_lp W=170n L=60n m=1
MNM6 net42 B net39 VSS nm1p2_lvt_lp W=170n L=60n m=1
MNM7 net39 A VSS VSS nm1p2_lvt_lp W=170n L=60n m=1
MPM4 net35 A VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM5 net35 B VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM6 net35 C VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM7 net35 D VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
XXI2 net35 VDD VSS Y / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND4X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND4X3H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MNM4 net35 D net45 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM5 net45 C net42 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM6 net42 B net39 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM7 net39 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM4 net35 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM5 net35 B VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM6 net35 C VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM7 net35 D VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI2 net35 VDD VSS Y / INV pl=6e-08 pw=5.7e-07 nl=6e-08 nw=4.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND4X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND4X4H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MNM0 net35 D net45 VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM1 net45 C net42 VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM2 net42 B net39 VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM3 net39 A VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MPM0 net35 A VDD VDD pm1p2_lvt_lp W=240n L=60n m=1
MPM1 net35 B VDD VDD pm1p2_lvt_lp W=240n L=60n m=1
MPM2 net35 C VDD VDD pm1p2_lvt_lp W=240n L=60n m=1
MPM3 net35 D VDD VDD pm1p2_lvt_lp W=240n L=60n m=1
XI0 net35 VDD VSS Y / INV pl=6e-08 pw=7.6e-07 nl=6e-08 nw=6e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AND4X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT AND4X6H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MNM0 net35 D net45 VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM1 net45 C net42 VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM2 net42 B net39 VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM3 net39 A VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MPM0 net35 A VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM1 net35 B VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM2 net35 C VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM3 net35 D VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
XI0 net35 VDD VSS Y / INV pl=6e-08 pw=11.4e-07 nl=6e-08 nw=9e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO211X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO211X0P5H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 net21 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net21 C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net5 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net21 A1 net5 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM3 net21 C0 net8 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net8 B0 net7 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net7 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net7 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net21 VDD VSS Y / INV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO211X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO211X0P7H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 net1 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net1 C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net7 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net1 A1 net7 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM3 net1 C0 net8 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net8 B0 net9 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net9 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net9 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net1 VDD VSS Y / INV pl=60n pw=222n nl=60n nw=174n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO211X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO211X1H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 net1 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net1 C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net7 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net1 A1 net7 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM3 net1 C0 net8 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net8 B0 net9 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net9 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net9 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net1 VDD VSS Y / INV pl=60n pw=270n nl=60n nw=210n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO211X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO211X1P4H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 net1 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net1 C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net7 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net1 A1 net7 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM3 net1 C0 net8 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net8 B0 net9 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net9 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net9 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net1 VDD VSS Y / INV pl=60n pw=314n nl=60n nw=246n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO211X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO211X2H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 net1 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net1 C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net7 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net1 A1 net7 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM3 net1 C0 net8 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net8 B0 net9 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net9 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net9 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net1 VDD VSS Y / INV pl=60n pw=380n nl=60n nw=300n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO211X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO211X3H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 net1 B0 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMNM2 net1 C0 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMNM1 net7 A0 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMNM0 net1 A1 net7 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMPM3 net1 C0 net8 VDD pm1p2_lvt_lp W=250n L=60n m=1
MMPM2 net8 B0 net9 VDD pm1p2_lvt_lp W=250n L=60n m=1
MMPM1 net9 A1 VDD VDD pm1p2_lvt_lp W=250n L=60n m=1
MMPM0 net9 A0 VDD VDD pm1p2_lvt_lp W=250n L=60n m=1
XXI1 net1 VDD VSS Y / INV pl=60n pw=570n nl=60n nw=450n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO211X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO211X4H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 net1 B0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM2 net1 C0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM1 net7 A0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM0 net1 A1 net7 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMPM3 net1 C0 net8 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM2 net8 B0 net9 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM1 net9 A1 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM0 net9 A0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
XXI1 net1 VDD VSS Y / INV pl=60n pw=760n nl=60n nw=600n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO211X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO211X6H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 net1 B0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM2 net1 C0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM1 net7 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM0 net1 A1 net7 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMPM3 net1 C0 net8 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM2 net8 B0 net9 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM1 net9 A1 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM0 net9 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
XXI1 net1 VDD VSS Y / INV pl=60n pw=1.14u nl=60n nw=0.9u
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO21X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO21X0P5H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMNM2 net17 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net25 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net17 A1 net25 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM2 net17 B0 net5 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net5 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net5 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net17 VDD VSS Y / INV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO21X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO21X0P7H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMNM2 net9 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net24 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net9 A1 net24 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM2 net9 B0 net19 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net19 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net19 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net9 VDD VSS Y / INV pl=60n pw=222n nl=60n nw=174n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO21X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO21X1H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMNM2 net9 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net24 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net9 A1 net24 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM2 net9 B0 net19 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net19 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net19 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net9 VDD VSS Y / INV pl=60n pw=270n nl=60n nw=210n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO21X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO21X1P4H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMNM2 net9 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net24 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net9 A1 net24 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM2 net9 B0 net19 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net19 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net19 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net9 VDD VSS Y / INV pl=60n pw=314n nl=60n nw=246n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO21X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO21X2H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMNM0 net8 A1 net23 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net23 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net8 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM0 net21 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net21 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net8 B0 net21 VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net8 VDD VSS Y / INV pl=60n pw=380n nl=60n nw=300n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO21X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO21X3H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMNM2 net9 B0 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMNM1 net24 A0 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMNM0 net9 A1 net24 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMPM2 net9 B0 net19 VDD pm1p2_lvt_lp W=250n L=60n m=1
MMPM1 net19 A1 VDD VDD pm1p2_lvt_lp W=250n L=60n m=1
MMPM0 net19 A0 VDD VDD pm1p2_lvt_lp W=250n L=60n m=1
XXI1 net9 VDD VSS Y / INV pl=60n pw=570n nl=60n nw=450n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO21X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO21X4H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMNM0 net42 A1 net55 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM1 net55 A0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM2 net42 B0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMPM0 net52 A0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM1 net52 A1 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM2 net42 B0 net52 VDD pm1p2_lvt_lp W=310n L=60n m=1
XXI1 net42 VDD VSS Y / INV pl=60n pw=760n nl=60n nw=600n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO21X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO21X6H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMNM2 net9 B0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM1 net24 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM0 net9 A1 net24 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMPM2 net9 B0 net19 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM1 net19 A1 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM0 net19 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
XXI1 net9 VDD VSS Y / INV pl=60n pw=1.14u nl=60n nw=0.9u
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO21X8H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO21X8H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMNM2 net9 B0 VSS VSS nm1p2_lvt_lp W=500n L=60n m=1
MMNM1 net24 A0 VSS VSS nm1p2_lvt_lp W=500n L=60n m=1
MMNM0 net9 A1 net24 VSS nm1p2_lvt_lp W=500n L=60n m=1
MMPM2 net9 B0 net19 VDD pm1p2_lvt_lp W=620n L=60n m=1
MMPM1 net19 A1 VDD VDD pm1p2_lvt_lp W=620n L=60n m=1
MMPM0 net19 A0 VDD VDD pm1p2_lvt_lp W=620n L=60n m=1
XXI1 net9 VDD VSS Y / INV pl=60n pw=1.52u nl=60n nw=1.2u
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO221X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO221X0P5H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MMNM4 net14 C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net31 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net14 B1 net31 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net39 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net14 A1 net39 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM4 net14 C0 net15 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net15 B1 net18 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net15 B0 net18 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net18 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net18 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net14 VDD VSS Y / INV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO221X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO221X0P7H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MMNM4 net1 C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net7 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net1 B1 net7 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net8 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net1 A1 net8 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM4 net1 C0 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net13 B1 net16 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net13 B0 net16 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net16 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net16 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net1 VDD VSS Y / INV pl=60n pw=222n nl=60n nw=174n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO221X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO221X1H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MMNM4 net1 C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net7 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net1 B1 net7 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net8 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net1 A1 net8 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM4 net1 C0 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net13 B1 net16 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net13 B0 net16 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net16 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net16 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net1 VDD VSS Y / INV pl=60n pw=270n nl=60n nw=210n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO221X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO221X1P4H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MMNM4 net1 C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net7 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net1 B1 net7 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net8 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net1 A1 net8 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM4 net1 C0 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net13 B1 net16 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net13 B0 net16 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net16 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net16 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net1 VDD VSS Y / INV pl=60n pw=314n nl=60n nw=246n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO221X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO221X2H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
XXI3 net52 VDD VSS Y / INV pl=60n pw=380n nl=60n nw=300n
MMPM3 net42 B1 net38 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM4 net52 C0 net42 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net42 B0 net38 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net38 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net38 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMNM0 net52 A1 net46 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net46 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM4 net52 C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net47 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net52 B1 net47 VSS nm1p2_lvt_lp W=150n L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO221X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO221X3H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MMNM4 net1 C0 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMNM3 net7 B0 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMNM2 net1 B1 net7 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMNM1 net8 A0 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMNM0 net1 A1 net8 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMPM4 net1 C0 net13 VDD pm1p2_lvt_lp W=250n L=60n m=1
MMPM3 net13 B1 net16 VDD pm1p2_lvt_lp W=250n L=60n m=1
MMPM2 net13 B0 net16 VDD pm1p2_lvt_lp W=250n L=60n m=1
MMPM1 net16 A1 VDD VDD pm1p2_lvt_lp W=250n L=60n m=1
MMPM0 net16 A0 VDD VDD pm1p2_lvt_lp W=250n L=60n m=1
XXI3 net1 VDD VSS Y / INV pl=60n pw=570n nl=60n nw=450n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO221X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO221X4H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MMNM4 net1 C0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM3 net7 B0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM2 net1 B1 net7 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM1 net8 A0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM0 net1 A1 net8 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMPM4 net1 C0 net13 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM3 net13 B1 net16 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM2 net13 B0 net16 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM1 net16 A1 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM0 net16 A0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
XXI3 net1 VDD VSS Y / INV pl=60n pw=760n nl=60n nw=600n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO222X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO222X0P5H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 net17 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM4 net44 A1 net17 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net32 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net44 B1 net32 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net48 C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net44 C1 net48 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM5 net44 C1 net19 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM4 net44 C0 net19 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net19 B1 net15 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net19 B0 net15 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net15 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net15 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net44 VDD VSS Y / INV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO222X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO222X0P7H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 net11 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM4 net1 A1 net11 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net10 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net1 B1 net10 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net6 C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net1 C1 net6 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM5 net1 C1 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM4 net1 C0 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net13 B1 net19 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net13 B0 net19 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net19 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net19 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net1 VDD VSS Y / INV pl=60n pw=222n nl=60n nw=174n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO222X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO222X1H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 net11 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM4 net1 A1 net11 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net10 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net1 B1 net10 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net6 C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net1 C1 net6 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM5 net1 C1 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM4 net1 C0 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net13 B1 net19 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net13 B0 net19 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net19 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net19 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net1 VDD VSS Y / INV pl=60n pw=270n nl=60n nw=210n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO222X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO222X1P4H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 net11 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM4 net1 A1 net11 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net10 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net1 B1 net10 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net6 C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net1 C1 net6 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM5 net1 C1 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM4 net1 C0 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net13 B1 net19 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net13 B0 net19 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net19 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net19 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net1 VDD VSS Y / INV pl=60n pw=314n nl=60n nw=246n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO222X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO222X2H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
XXI1 net4 VDD VSS Y / INV pl=60n pw=380n nl=60n nw=300n
MMPM4 net4 C0 net48 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM5 net4 C1 net48 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net48 B1 net42 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net48 B0 net42 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net42 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net42 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMNM0 net4 C1 net57 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net57 C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net4 B1 net53 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net53 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM4 net4 A1 net52 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM5 net52 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO222X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO222X3H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 net11 A0 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMNM4 net1 A1 net11 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMNM3 net10 B0 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMNM2 net1 B1 net10 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMNM1 net6 C0 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMNM0 net1 C1 net6 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMPM5 net1 C1 net13 VDD pm1p2_lvt_lp W=250n L=60n m=1
MMPM4 net1 C0 net13 VDD pm1p2_lvt_lp W=250n L=60n m=1
MMPM3 net13 B1 net19 VDD pm1p2_lvt_lp W=250n L=60n m=1
MMPM2 net13 B0 net19 VDD pm1p2_lvt_lp W=250n L=60n m=1
MMPM1 net19 A1 VDD VDD pm1p2_lvt_lp W=250n L=60n m=1
MMPM0 net19 A0 VDD VDD pm1p2_lvt_lp W=250n L=60n m=1
XXI1 net1 VDD VSS Y / INV pl=60n pw=570n nl=60n nw=450n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO222X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO222X4H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 net11 A0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM4 net1 A1 net11 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM3 net10 B0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM2 net1 B1 net10 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM1 net6 C0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM0 net1 C1 net6 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMPM5 net1 C1 net13 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM4 net1 C0 net13 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM3 net13 B1 net19 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM2 net13 B0 net19 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM1 net19 A1 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM0 net19 A0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
XXI1 net1 VDD VSS Y / INV pl=60n pw=760n nl=60n nw=600n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO22X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO22X0P5H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MMNM3 net9 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net13 A1 net9 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net8 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net13 B1 net8 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM3 net13 B1 net17 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net17 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net13 B0 net17 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net17 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net13 VDD VSS Y / INV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO22X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO22X0P7H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MMNM3 net13 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net1 A1 net13 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net14 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net1 B1 net14 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM3 net1 B1 net8 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net8 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net1 B0 net8 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net8 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net1 VDD VSS Y / INV pl=60n pw=222n nl=60n nw=174n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO22X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO22X1H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MMNM3 net13 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net1 A1 net13 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net14 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net1 B1 net14 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM3 net1 B1 net8 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net8 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net1 B0 net8 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net8 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net1 VDD VSS Y / INV pl=60n pw=270n nl=60n nw=210n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO22X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO22X1P4H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MMNM3 net13 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net1 A1 net13 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net14 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net1 B1 net14 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM3 net1 B1 net8 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net8 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net1 B0 net8 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net8 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net1 VDD VSS Y / INV pl=60n pw=314n nl=60n nw=246n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO22X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO22X2H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MMNM0 net42 B1 net30 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net30 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net42 A1 net31 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net31 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM0 net35 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net42 B0 net35 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net35 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net42 B1 net35 VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net42 VDD VSS Y / INV pl=60n pw=380n nl=60n nw=300n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO22X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO22X3H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MMNM3 net13 A0 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMNM2 net1 A1 net13 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMNM1 net14 B0 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMNM0 net1 B1 net14 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMPM3 net1 B1 net8 VDD pm1p2_lvt_lp W=250n L=60n m=1
MMPM2 net8 A1 VDD VDD pm1p2_lvt_lp W=250n L=60n m=1
MMPM1 net1 B0 net8 VDD pm1p2_lvt_lp W=250n L=60n m=1
MMPM0 net8 A0 VDD VDD pm1p2_lvt_lp W=250n L=60n m=1
XXI1 net1 VDD VSS Y / INV pl=60n pw=570n nl=60n nw=450n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO22X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO22X4H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
XXI1 net1 VDD VSS Y / INV pl=60n pw=760n nl=60n nw=600n
MMPM1 net1 B0 net8 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM0 net8 A0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM2 net8 A1 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM3 net1 B1 net8 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMNM3 net13 A0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM2 net1 A1 net13 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM0 net1 B1 net14 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM1 net14 B0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO22X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO22X6H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MMNM3 net13 A0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM2 net1 A1 net13 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM1 net14 B0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM0 net1 B1 net14 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMPM3 net1 B1 net8 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM2 net8 A1 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM1 net1 B0 net8 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM0 net8 A0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
XXI1 net1 VDD VSS Y / INV pl=60n pw=1.14u nl=60n nw=900n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO31X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO31X0P5H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMNM3 net36 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net28 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net13 A1 net28 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net36 A2 net13 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM3 net36 B0 net8 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net8 A2 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net8 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net8 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net36 VDD VSS Y / INV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO31X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO31X0P7H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMNM3 net1 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net11 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net10 A1 net11 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net1 A2 net10 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM3 net1 B0 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net13 A2 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net13 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net1 VDD VSS Y / INV pl=60n pw=222n nl=60n nw=174n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO31X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO31X1H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMNM3 net1 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net11 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net10 A1 net11 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net1 A2 net10 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM3 net1 B0 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net13 A2 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net13 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net1 VDD VSS Y / INV pl=60n pw=270n nl=60n nw=210n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO31X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO31X1P4H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMNM3 net1 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net11 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net10 A1 net11 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net1 A2 net10 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM3 net1 B0 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net13 A2 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net13 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net1 VDD VSS Y / INV pl=60n pw=314n nl=60n nw=246n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO31X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO31X2H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
XXI3 net35 VDD VSS Y / INV pl=60n pw=380n nl=60n nw=300n
MMPM2 net42 A2 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net35 B0 net42 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net42 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net42 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMNM0 net35 A2 net34 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net34 A1 net33 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net35 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net33 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO31X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO31X3H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMNM3 net1 B0 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMNM2 net11 A0 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMNM1 net10 A1 net11 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMNM0 net1 A2 net10 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMPM3 net1 B0 net13 VDD pm1p2_lvt_lp W=250n L=60n m=1
MMPM2 net13 A2 VDD VDD pm1p2_lvt_lp W=250n L=60n m=1
MMPM1 net13 A1 VDD VDD pm1p2_lvt_lp W=250n L=60n m=1
MMPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=250n L=60n m=1
XXI3 net1 VDD VSS Y / INV pl=60n pw=570n nl=60n nw=450n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AO31X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AO31X4H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMNM3 net1 B0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM2 net11 A0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM1 net10 A1 net11 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM0 net1 A2 net10 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMPM3 net1 B0 net13 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM2 net13 A2 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM1 net13 A1 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
XXI3 net1 VDD VSS Y / INV pl=60n pw=760n nl=60n nw=600n
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOA211X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOA211X0P5H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM5 net6 B0 net19 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM1 net19 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM2 net19 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM0 net6 C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM14 Y net6 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM4 net16 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM6 net16 A0 net30 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM7 net6 C0 net16 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM3 net30 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM13 Y net6 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOA211X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOA211X0P7H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM5 net6 B0 net10 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM1 net10 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM2 net10 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM0 net6 C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM14 Y net6 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMM4 net26 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM6 net26 A0 net38 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM7 net6 C0 net26 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM3 net38 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM13 Y net6 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOA211X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOA211X1H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM5 net6 B0 net10 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM1 net10 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM2 net10 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM0 net6 C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM14 Y net6 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMM4 net26 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM6 net26 A0 net38 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM7 net6 C0 net26 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM3 net38 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM13 Y net6 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOA211X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOA211X1P4H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM5 net6 B0 net10 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM1 net10 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM2 net10 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM0 net6 C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM14 Y net6 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMM4 net26 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM6 net26 A0 net38 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM7 net6 C0 net26 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM3 net38 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM13 Y net6 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOA211X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOA211X2H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM5 net6 B0 net10 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM1 net10 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM2 net10 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM0 net6 C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM14 Y net6 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMM4 net26 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM6 net26 A0 net38 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM7 net6 C0 net26 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM3 net38 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM13 Y net6 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOA211X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOA211X3H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM5 net6 B0 net10 VDD pm1p2_lvt_lp W=250n L=60n m=1
MMM1 net10 A0 VDD VDD pm1p2_lvt_lp W=250n L=60n m=1
MMM2 net10 A1 VDD VDD pm1p2_lvt_lp W=250n L=60n m=1
MMM0 net6 C0 VDD VDD pm1p2_lvt_lp W=250n L=60n m=1
MMM14 Y net6 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMM4 net26 B0 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMM6 net26 A0 net38 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMM7 net6 C0 net26 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMM3 net38 A1 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMM13 Y net6 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOA211X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOA211X4H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM5 net6 B0 net10 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMM1 net10 A0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MMM2 net10 A1 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MMM0 net6 C0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MMM14 Y net6 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMM4 net26 B0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMM6 net26 A0 net38 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMM7 net6 C0 net26 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMM3 net38 A1 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMM13 Y net6 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOAI211X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOAI211X0P5H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM3 net21 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM7 Y C0 net19 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM6 net19 A0 net21 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM4 net19 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM0 Y C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM2 net8 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM1 net8 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM5 Y B0 net8 VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOAI211X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOAI211X0P7H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM3 net21 A1 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMM7 Y C0 net19 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMM6 net19 A0 net21 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMM4 net19 B0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMM0 Y C0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMM2 net8 A1 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMM1 net8 A0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMM5 Y B0 net8 VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOAI211X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOAI211X1H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM3 net21 A1 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMM7 Y C0 net19 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMM6 net19 A0 net21 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMM4 net19 B0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMM0 Y C0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMM2 net8 A1 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMM1 net8 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMM5 Y B0 net8 VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOAI211X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOAI211X1P4H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM3 net21 A1 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMM7 Y C0 net19 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMM6 net19 A0 net21 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMM4 net19 B0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMM0 Y C0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMM2 net8 A1 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMM1 net8 A0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMM5 Y B0 net8 VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOAI211X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOAI211X2H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM3 net21 A1 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMM7 Y C0 net19 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMM6 net19 A0 net21 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMM4 net19 B0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMM0 Y C0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMM2 net8 A1 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMM1 net8 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMM5 Y B0 net8 VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOAI211X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOAI211X3H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM3 net21 A1 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMM7 Y C0 net19 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMM6 net19 A0 net21 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMM4 net19 B0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMM0 Y C0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMM2 net8 A1 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMM1 net8 A0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMM5 Y B0 net8 VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOAI211X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOAI211X4H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM3 net21 A1 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMM7 Y C0 net19 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMM6 net19 A0 net21 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMM4 net19 B0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMM0 Y C0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMM2 net8 A1 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMM1 net8 A0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMM5 Y B0 net8 VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI211X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI211X0P5H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMN5 Y B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net13 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 Y A1 net13 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 Y C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP3 Y B0 net8 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP2 net8 C0 net039 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 net039 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP0 net039 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI211X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI211X0P7H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMN5 Y B0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN4 net7 A0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN1 Y A1 net7 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN0 Y C0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMP3 Y B0 net8 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP2 net8 C0 net9 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP1 net9 A1 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP0 net9 A0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI211X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI211X1H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMN5 Y B0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN4 net7 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN1 Y A1 net7 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN0 Y C0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMP3 Y B0 net8 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP2 net8 C0 net9 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP1 net9 A1 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP0 net9 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI211X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI211X1P4H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMN5 Y B0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN4 net7 A0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN1 Y A1 net7 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN0 Y C0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMP3 Y B0 net8 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP2 net8 C0 net9 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP1 net9 A1 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP0 net9 A0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI211X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI211X2H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMN0 Y C0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN1 Y A1 net34 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN4 net34 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN5 Y B0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP0 net31 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP1 net31 A1 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP2 net33 C0 net31 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP3 Y B0 net33 VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI211X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI211X3H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMN5 Y B0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN4 net7 A0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN1 Y A1 net7 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN0 Y C0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMP3 Y B0 net8 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP2 net8 C0 net9 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP1 net9 A1 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP0 net9 A0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI211X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI211X4H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMP1 net9 A1 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP0 net9 A0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP2 net8 C0 net9 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP3 Y B0 net8 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMN5 Y B0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN4 net7 A0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN1 Y A1 net7 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN0 Y C0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI211X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI211X6H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMN5 Y B0 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN4 net7 A0 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN1 Y A1 net7 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN0 Y C0 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMP3 Y B0 net8 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP2 net8 C0 net9 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP1 net9 A1 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP0 net9 A0 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI21BX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI21BX0P5H7L A0 A1 B0N VDD VSS Y
*.PININFO A0:I A1:I B0N:I Y:O VDD:B VSS:B
MMNM2 Y net066 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net8 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 Y A1 net8 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM2 Y net066 net5 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net5 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net5 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI4 B0N VDD VSS net066 / INV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI21BX0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI21BX0P7H7L A0 A1 B0N VDD VSS Y
*.PININFO A0:I A1:I B0N:I Y:O VDD:B VSS:B
MMNM2 Y net066 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM1 net9 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 Y A1 net9 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM2 Y net066 net8 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM1 net8 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net8 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI4 B0N VDD VSS net066 / INV pl=60n pw=222n nl=60n nw=174n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI21BX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI21BX1H7L A0 A1 B0N VDD VSS Y
*.PININFO A0:I A1:I B0N:I Y:O VDD:B VSS:B
MMNM2 Y net066 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM1 net9 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 Y A1 net9 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM2 Y net066 net8 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM1 net8 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net8 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI4 B0N VDD VSS net066 / INV pl=60n pw=270n nl=60n nw=210n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI21BX1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI21BX1P4H7L A0 A1 B0N VDD VSS Y
*.PININFO A0:I A1:I B0N:I Y:O VDD:B VSS:B
MMNM2 Y net066 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM1 net9 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 Y A1 net9 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM2 Y net066 net8 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM1 net8 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net8 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI4 B0N VDD VSS net066 / INV pl=60n pw=314n nl=60n nw=246n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI21BX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI21BX2H7L A0 A1 B0N VDD VSS Y
*.PININFO A0:I A1:I B0N:I Y:O VDD:B VSS:B
MMNM2 Y net066 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM1 net9 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 Y A1 net9 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM2 Y net066 net8 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM1 net8 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net8 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI4 B0N VDD VSS net066 / INV pl=60n pw=380n nl=60n nw=300n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI21BX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI21BX3H7L A0 A1 B0N VDD VSS Y
*.PININFO A0:I A1:I B0N:I Y:O VDD:B VSS:B
MMNM2 Y net066 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM1 net9 A0 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMNM0 Y A1 net9 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMPM2 Y net066 net8 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM1 net8 A1 VDD VDD pm1p2_lvt_lp W=250n L=60n m=1
MMPM0 net8 A0 VDD VDD pm1p2_lvt_lp W=250n L=60n m=1
XXI4 B0N VDD VSS net066 / INV pl=60n pw=570n nl=60n nw=450n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI21BX4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI21BX4H7L A0 A1 B0N VDD VSS Y
*.PININFO A0:I A1:I B0N:I Y:O VDD:B VSS:B
MMNM2 Y net066 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM1 net9 A0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM0 Y A1 net9 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMPM2 Y net066 net8 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM1 net8 A1 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM0 net8 A0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
XXI4 B0N VDD VSS net066 / INV pl=60n pw=760n nl=60n nw=600n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI21BX6H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI21BX6H7L A0 A1 B0N VDD VSS Y
*.PININFO A0:I A1:I B0N:I Y:O VDD:B VSS:B
MMNM2 Y net066 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMNM1 net9 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM0 Y A1 net9 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMPM2 Y net066 net8 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMPM1 net8 A1 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM0 net8 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
XXI4 B0N VDD VSS net066 / INV pl=60n pw=1.14u nl=60n nw=0.9u
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI21X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI21X0P5H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMN4 net5 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 Y A1 net5 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 Y B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP2 Y B0 net8 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 net8 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP0 net8 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI21X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI21X0P7H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMP1 net31 A1 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP2 Y B0 net31 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP0 net31 A0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMN0 Y B0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN1 Y A1 net33 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN4 net33 A0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI21X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI21X1H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMP1 net31 A1 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP2 Y B0 net31 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP0 net31 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMN0 Y B0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN1 Y A1 net33 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN4 net33 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI21X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI21X1P4H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMP1 net31 A1 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP2 Y B0 net31 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP0 net31 A0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMN0 Y B0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN1 Y A1 net33 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN4 net33 A0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI21X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI21X2H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMN4 net60 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN1 Y A1 net60 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN0 Y B0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP2 Y B0 net59 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP1 net59 A1 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP0 net59 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI21X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI21X3H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMP1 net31 A1 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP2 Y B0 net31 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP0 net31 A0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMN0 Y B0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN1 Y A1 net33 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN4 net33 A0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI21X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI21X4H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMN4 net60 A0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN1 Y A1 net60 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN0 Y B0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMP2 Y B0 net59 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP1 net59 A1 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP0 net59 A0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI21X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI21X6H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMP1 net31 A1 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP2 Y B0 net31 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP0 net31 A0 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMN0 Y B0 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN1 Y A1 net33 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN4 net33 A0 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI21X8H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI21X8H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMP1 net31 A1 VDD VDD pm1p2_lvt_lp W=1.52u L=60n m=1
MMP2 Y B0 net31 VDD pm1p2_lvt_lp W=1.52u L=60n m=1
MMP0 net31 A0 VDD VDD pm1p2_lvt_lp W=1.52u L=60n m=1
MMN0 Y B0 VSS VSS nm1p2_lvt_lp W=1.2u L=60n m=1
MMN1 Y A1 net33 VSS nm1p2_lvt_lp W=1.2u L=60n m=1
MMN4 net33 A0 VSS VSS nm1p2_lvt_lp W=1.2u L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI221X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI221X0P5H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MMNM4 Y C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net31 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 Y B1 net31 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net1 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 Y A1 net1 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM4 Y C0 net7 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net7 B1 net5 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net7 B0 net5 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net5 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net5 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI221X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI221X0P7H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MMNM4 Y C0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM3 net16 B0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM2 Y B1 net16 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM1 net17 A0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM0 Y A1 net17 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMPM4 Y C0 net1 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM3 net1 B1 net8 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM2 net1 B0 net8 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM1 net8 A1 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM0 net8 A0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI221X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI221X1H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MMNM4 Y C0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM3 net16 B0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM2 Y B1 net16 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM1 net17 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM0 Y A1 net17 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMPM4 Y C0 net1 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM3 net1 B1 net8 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM2 net1 B0 net8 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM1 net8 A1 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM0 net8 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI221X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI221X1P4H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MMNM4 Y C0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM3 net16 B0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM2 Y B1 net16 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM1 net17 A0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM0 Y A1 net17 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMPM4 Y C0 net1 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM3 net1 B1 net8 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM2 net1 B0 net8 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM1 net8 A1 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM0 net8 A0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI221X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI221X2H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MMPM3 net48 B1 net42 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM4 Y C0 net48 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM2 net48 B0 net42 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM0 net42 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM1 net42 A1 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMNM0 Y A1 net34 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM1 net34 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM2 Y B1 net35 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM3 net35 B0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM4 Y C0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI221X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI221X3H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MMNM4 Y C0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM3 net16 B0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM2 Y B1 net16 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM1 net17 A0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM0 Y A1 net17 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMPM4 Y C0 net1 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM3 net1 B1 net8 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM2 net1 B0 net8 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM1 net8 A1 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM0 net8 A0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI221X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI221X4H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MMNM4 Y C0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM3 net16 B0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM2 Y B1 net16 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM1 net17 A0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM0 Y A1 net17 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMPM4 Y C0 net1 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM3 net1 B1 net8 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM2 net1 B0 net8 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM1 net8 A1 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM0 net8 A0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI222X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI222X0P5H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 net40 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM4 Y A1 net40 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net32 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 Y B1 net32 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net48 C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 Y C1 net48 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM5 Y C1 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM4 Y C0 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net13 B1 net15 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net13 B0 net15 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net15 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net15 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI222X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI222X0P7H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 net14 A0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM4 Y A1 net14 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM3 net52 B0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM2 Y B1 net52 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM1 net51 C0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM0 Y C1 net51 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMPM5 Y C1 net54 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM4 Y C0 net54 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM3 net54 B1 net45 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM2 net54 B0 net45 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM1 net45 A1 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM0 net45 A0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI222X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI222X1H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 net14 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM4 Y A1 net14 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM3 net52 B0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM2 Y B1 net52 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM1 net51 C0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM0 Y C1 net51 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMPM5 Y C1 net54 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM4 Y C0 net54 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM3 net54 B1 net45 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM2 net54 B0 net45 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM1 net45 A1 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM0 net45 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI222X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI222X1P4H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 net14 A0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM4 Y A1 net14 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM3 net52 B0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM2 Y B1 net52 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM1 net51 C0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM0 Y C1 net51 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMPM5 Y C1 net54 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM4 Y C0 net54 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM3 net54 B1 net45 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM2 net54 B0 net45 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM1 net45 A1 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM0 net45 A0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI222X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI222X2H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMPM4 Y C0 net1 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM5 Y C1 net1 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM3 net1 B1 net13 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM1 net13 A1 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM2 net1 B0 net13 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMNM0 Y C1 net9 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM1 net9 C0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM2 Y B1 net8 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM3 net8 B0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM4 Y A1 net46 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM5 net46 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI222X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI222X3H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 net14 A0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM4 Y A1 net14 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM3 net52 B0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM2 Y B1 net52 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM1 net51 C0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM0 Y C1 net51 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMPM5 Y C1 net54 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM4 Y C0 net54 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM3 net54 B1 net45 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM2 net54 B0 net45 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM1 net45 A1 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM0 net45 A0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI222X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI222X4H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 net14 A0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM4 Y A1 net14 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM3 net52 B0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM2 Y B1 net52 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM1 net51 C0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM0 Y C1 net51 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMPM5 Y C1 net54 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM4 Y C0 net54 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM3 net54 B1 net45 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM2 net54 B0 net45 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM1 net45 A1 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM0 net45 A0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI22X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI22X0P5H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MMN5 net8 B1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net9 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 Y A1 net9 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 Y B0 net8 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP3 Y B1 net051 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP2 Y B0 net051 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 net051 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP0 net051 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI22X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI22X0P7H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MMN5 net14 B1 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN4 net13 A0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN1 Y A1 net13 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN0 Y B0 net14 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMP3 Y B1 net8 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP2 Y B0 net8 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP1 net8 A1 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP0 net8 A0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI22X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI22X1H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MMN5 net14 B1 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN4 net13 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN1 Y A1 net13 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN0 Y B0 net14 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMP3 Y B1 net8 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP2 Y B0 net8 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP1 net8 A1 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP0 net8 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI22X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI22X1P4H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MMN5 net14 B1 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN4 net13 A0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN1 Y A1 net13 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN0 Y B0 net14 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMP3 Y B1 net8 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP2 Y B0 net8 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP1 net8 A1 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP0 net8 A0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI22X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI22X2H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MMP2 Y B0 net31 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP3 Y B1 net31 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP1 net31 A1 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP0 net31 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMN0 Y B0 net27 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN1 Y A1 net28 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN4 net28 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN5 net27 B1 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI22X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI22X3H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MMN5 net14 B1 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN4 net13 A0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN1 Y A1 net13 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN0 Y B0 net14 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMP3 Y B1 net8 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP2 Y B0 net8 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP1 net8 A1 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP0 net8 A0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI22X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI22X4H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MMN5 net14 B1 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN4 net13 A0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN1 Y A1 net13 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN0 Y B0 net14 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMP3 Y B1 net8 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP2 Y B0 net8 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP1 net8 A1 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP0 net8 A0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI22X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI22X6H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MMN5 net14 B1 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN4 net13 A0 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN1 Y A1 net13 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN0 Y B0 net14 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMP3 Y B1 net8 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP2 Y B0 net8 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP1 net8 A1 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP0 net8 A0 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2BB1X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2BB1X0P5H7L A0N A1N B0 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I Y:O VDD:B VSS:B
MMN5 net8 A0N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 Y B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN7 Y net8 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN6 net8 A1N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP4 net8 A1N net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP3 net13 A0N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP2 Y B0 net12 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 net12 net8 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2BB1X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2BB1X0P7H7L A0N A1N B0 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I Y:O VDD:B VSS:B
MMN6 net42 A1N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN7 Y net42 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN4 Y B0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN5 net42 A0N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP1 net40 net42 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP2 Y B0 net40 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP3 net39 A0N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP4 net42 A1N net39 VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2BB1X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2BB1X1H7L A0N A1N B0 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I Y:O VDD:B VSS:B
MMN6 net42 A1N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN7 Y net42 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN4 Y B0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN5 net42 A0N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP1 net40 net42 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP2 Y B0 net40 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP3 net39 A0N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP4 net42 A1N net39 VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2BB1X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2BB1X1P4H7L A0N A1N B0 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I Y:O VDD:B VSS:B
MMN6 net42 A1N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN7 Y net42 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN4 Y B0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN5 net42 A0N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP1 net40 net42 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP2 Y B0 net40 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP3 net39 A0N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP4 net42 A1N net39 VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2BB1X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2BB1X2H7L A0N A1N B0 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I Y:O VDD:B VSS:B
MMN6 net54 A1N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN7 Y net54 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN4 Y B0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN5 net54 A0N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP1 net56 net54 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP2 Y B0 net56 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP3 net57 A0N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP4 net54 A1N net57 VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2BB1X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2BB1X3H7L A0N A1N B0 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I Y:O VDD:B VSS:B
MMN6 net42 A1N VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN7 Y net42 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN4 Y B0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN5 net42 A0N VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMP1 net40 net42 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP2 Y B0 net40 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP3 net39 A0N VDD VDD pm1p2_lvt_lp W=250n L=60n m=1
MMP4 net42 A1N net39 VDD pm1p2_lvt_lp W=250n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2BB1X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2BB1X4H7L A0N A1N B0 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I Y:O VDD:B VSS:B
MMP4 net75 A1N net73 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMP3 net73 A0N VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MMP2 Y B0 net74 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP1 net74 net75 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMN5 net75 A0N VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMN4 Y B0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN7 Y net75 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN6 net75 A1N VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2BB1X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2BB1X6H7L A0N A1N B0 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I Y:O VDD:B VSS:B
MMN6 net42 A1N VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN7 Y net42 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN4 Y B0 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN5 net42 A0N VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP1 net40 net42 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP2 Y B0 net40 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP3 net39 A0N VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP4 net42 A1N net39 VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2BB2X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2BB2X0P5H7L A0N A1N B0 B1 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I B1:I Y:O VDD:B VSS:B
MMN5 net8 A1N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN6 Y net8 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net15 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 Y B1 net15 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 net8 A0N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP5 Y net8 net053 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP4 net053 B1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP3 net8 A1N net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP2 net053 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP0 net13 A0N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2BB2X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2BB2X0P7H7L A0N A1N B0 B1 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I B1:I Y:O VDD:B VSS:B
MMN5 net8 A1N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN6 Y net8 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN4 net10 B0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN1 Y B1 net10 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN0 net8 A0N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP5 Y net8 net13 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP4 net13 B1 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP3 net8 A1N net15 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP2 net13 B0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP0 net15 A0N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2BB2X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2BB2X1H7L A0N A1N B0 B1 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I B1:I Y:O VDD:B VSS:B
MMN5 net8 A1N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN6 Y net8 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN4 net10 B0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN1 Y B1 net10 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN0 net8 A0N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP5 Y net8 net13 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP4 net13 B1 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP3 net8 A1N net15 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP2 net13 B0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP0 net15 A0N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2BB2X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2BB2X1P4H7L A0N A1N B0 B1 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I B1:I Y:O VDD:B VSS:B
MMN5 net8 A1N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN6 Y net8 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN4 net10 B0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN1 Y B1 net10 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN0 net8 A0N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP5 Y net8 net13 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP4 net13 B1 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP3 net8 A1N net15 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP2 net13 B0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP0 net15 A0N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2BB2X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2BB2X2H7L A0N A1N B0 B1 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I B1:I Y:O VDD:B VSS:B
MMN5 net8 A1N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN6 Y net8 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN4 net10 B0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN1 Y B1 net10 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN0 net8 A0N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP5 Y net8 net13 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP4 net13 B1 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP3 net8 A1N net15 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP2 net13 B0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP0 net15 A0N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2BB2X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2BB2X3H7L A0N A1N B0 B1 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I B1:I Y:O VDD:B VSS:B
MMN5 net8 A1N VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN6 Y net8 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN4 net10 B0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN1 Y B1 net10 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN0 net8 A0N VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMP5 Y net8 net13 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP4 net13 B1 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP3 net8 A1N net15 VDD pm1p2_lvt_lp W=250n L=60n m=1
MMP2 net13 B0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP0 net15 A0N VDD VDD pm1p2_lvt_lp W=250n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2BB2X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2BB2X4H7L A0N A1N B0 B1 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I B1:I Y:O VDD:B VSS:B
MMN5 net8 A1N VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMN6 Y net8 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN4 net10 B0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN1 Y B1 net10 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN0 net8 A0N VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMP5 Y net8 net13 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP4 net13 B1 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP3 net8 A1N net15 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMP2 net13 B0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP0 net15 A0N VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2BB2X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2BB2X6H7L A0N A1N B0 B1 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I B1:I Y:O VDD:B VSS:B
MMN5 net8 A1N VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN6 Y net8 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN4 net10 B0 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN1 Y B1 net10 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN0 net8 A0N VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP5 Y net8 net13 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP4 net13 B1 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP3 net8 A1N net15 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP2 net13 B0 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP0 net15 A0N VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2XB1X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2XB1X0P5H7L A0 A1N B0 VDD VSS Y
*.PININFO A0:I A1N:I B0:I Y:O VDD:B VSS:B
MMNM3 net15 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 Y net6 net15 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 Y B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM2 Y B0 net14 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net14 net6 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net14 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 A1N VDD VSS net6 / INV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2XB1X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2XB1X0P7H7L A0 A1N B0 VDD VSS Y
*.PININFO A0:I A1N:I B0:I Y:O VDD:B VSS:B
MMNM3 net15 A0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM2 Y net6 net15 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM0 Y B0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMPM2 Y B0 net1 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM1 net1 net6 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM0 net1 A0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
XXI3 A1N VDD VSS net6 / INV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2XB1X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2XB1X1H7L A0 A1N B0 VDD VSS Y
*.PININFO A0:I A1N:I B0:I Y:O VDD:B VSS:B
MMNM3 net15 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM2 Y net6 net15 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM0 Y B0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMPM2 Y B0 net8 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM1 net8 net6 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM0 net8 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
XXI3 A1N VDD VSS net6 / INV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2XB1X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2XB1X1P4H7L A0 A1N B0 VDD VSS Y
*.PININFO A0:I A1N:I B0:I Y:O VDD:B VSS:B
MMNM3 net15 A0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM2 Y net6 net15 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM0 Y B0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMPM2 Y B0 net1 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM1 net1 net6 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM0 net1 A0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
XXI3 A1N VDD VSS net6 / INV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2XB1X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2XB1X2H7L A0 A1N B0 VDD VSS Y
*.PININFO A0:I A1N:I B0:I Y:O VDD:B VSS:B
MMNM3 net15 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM2 Y net6 net15 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM0 Y B0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMPM2 Y B0 net8 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM1 net8 net6 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM0 net8 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
XXI3 A1N VDD VSS net6 / INV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2XB1X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2XB1X3H7L A0 A1N B0 VDD VSS Y
*.PININFO A0:I A1N:I B0:I Y:O VDD:B VSS:B
MMNM3 net15 A0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM2 Y net6 net15 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM0 Y B0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMPM2 Y B0 net1 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM1 net1 net6 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM0 net1 A0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
XXI3 A1N VDD VSS net6 / INV pl=60n pw=250n nl=60n nw=200n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2XB1X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2XB1X4H7L A0 A1N B0 VDD VSS Y
*.PININFO A0:I A1N:I B0:I Y:O VDD:B VSS:B
MMNM3 net15 A0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM2 Y net6 net15 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM0 Y B0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMPM2 Y B0 net8 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM1 net8 net6 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM0 net8 A0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
XXI3 A1N VDD VSS net6 / INV pl=60n pw=310n nl=60n nw=250n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI2XB1X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI2XB1X6H7L A0 A1N B0 VDD VSS Y
*.PININFO A0:I A1N:I B0:I Y:O VDD:B VSS:B
MMNM3 net15 A0 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMNM2 Y net6 net15 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMNM0 Y B0 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMPM2 Y B0 net1 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMPM1 net1 net6 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMPM0 net1 A0 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
XXI3 A1N VDD VSS net6 / INV pl=60n pw=380n nl=60n nw=300n
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI31X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI31X0P5H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMN5 net37 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net12 A1 net37 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 Y A2 net12 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 Y B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP2 Y B0 net8 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP3 net8 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 net8 A2 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP0 net8 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI31X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI31X0P7H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMN5 net6 A0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN4 net5 A1 net6 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN1 Y A2 net5 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN0 Y B0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMP2 Y B0 net8 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP3 net8 A1 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP1 net8 A2 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP0 net8 A0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI31X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI31X1H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMN5 net6 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN4 net5 A1 net6 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN1 Y A2 net5 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN0 Y B0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMP2 Y B0 net8 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP3 net8 A1 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP1 net8 A2 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP0 net8 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI31X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI31X1P4H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMN5 net6 A0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN4 net5 A1 net6 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN1 Y A2 net5 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN0 Y B0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMP2 Y B0 net8 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP3 net8 A1 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP1 net8 A2 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP0 net8 A0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI31X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI31X2H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMP3 net31 A1 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP2 Y B0 net31 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP1 net31 A2 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP0 net31 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMN0 Y B0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN1 Y A2 net36 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN4 net36 A1 net35 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN5 net35 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI31X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI31X3H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMN5 net6 A0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN4 net5 A1 net6 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN1 Y A2 net5 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN0 Y B0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMP2 Y B0 net8 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP3 net8 A1 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP1 net8 A2 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP0 net8 A0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI31X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI31X4H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMN5 net6 A0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN4 net5 A1 net6 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN1 Y A2 net5 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN0 Y B0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMP2 Y B0 net8 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP3 net8 A1 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP1 net8 A2 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP0 net8 A0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI32X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI32X0P5H7L A0 A1 A2 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I Y:O VDD:B VSS:B
MMN5 net37 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN6 net45 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net12 A1 net37 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 Y A2 net12 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 Y B1 net45 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP4 Y B0 net19 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP3 net19 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP2 Y B1 net19 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 net19 A2 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP0 net19 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI32X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI32X0P7H7L A0 A1 A2 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I Y:O VDD:B VSS:B
MMN5 net17 A0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN6 net15 B0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN4 net16 A1 net17 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN1 Y A2 net16 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN0 Y B1 net15 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMP4 Y B0 net8 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP3 net8 A1 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP2 Y B1 net8 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP1 net8 A2 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP0 net8 A0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI32X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI32X1H7L A0 A1 A2 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I Y:O VDD:B VSS:B
MMN5 net17 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN6 net15 B0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN4 net16 A1 net17 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN1 Y A2 net16 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN0 Y B1 net15 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMP4 Y B0 net8 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP3 net8 A1 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP2 Y B1 net8 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP1 net8 A2 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP0 net8 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI32X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI32X1P4H7L A0 A1 A2 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I Y:O VDD:B VSS:B
MMN5 net17 A0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN6 net15 B0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN4 net16 A1 net17 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN1 Y A2 net16 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN0 Y B1 net15 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMP4 Y B0 net8 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP3 net8 A1 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP2 Y B1 net8 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP1 net8 A2 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP0 net8 A0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI32X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI32X2H7L A0 A1 A2 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I Y:O VDD:B VSS:B
MMP3 net42 A1 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP4 Y B0 net42 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP2 Y B1 net42 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP0 net42 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP1 net42 A2 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMN0 Y B1 net36 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN1 Y A2 net35 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN4 net35 A1 net34 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN6 net36 B0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN5 net34 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI32X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI32X3H7L A0 A1 A2 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I Y:O VDD:B VSS:B
MMN5 net17 A0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN6 net15 B0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN4 net16 A1 net17 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN1 Y A2 net16 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN0 Y B1 net15 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMP4 Y B0 net8 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP3 net8 A1 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP2 Y B1 net8 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP1 net8 A2 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP0 net8 A0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI32X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI32X4H7L A0 A1 A2 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I Y:O VDD:B VSS:B
MMN5 net17 A0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN6 net15 B0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN4 net16 A1 net17 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN1 Y A2 net16 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN0 Y B1 net15 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMP4 Y B0 net8 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP3 net8 A1 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP2 Y B1 net8 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP1 net8 A2 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP0 net8 A0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI33X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI33X0P5H7L A0 A1 A2 B0 B1 B2 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I B2:I Y:O VDD:B VSS:B
MMNM5 Y A2 net40 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM4 Y B2 net44 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net40 A1 net48 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net44 B1 net13 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net48 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net13 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM5 Y B1 net31 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM4 net31 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net31 A2 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net31 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 Y B2 net31 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 Y B0 net31 VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI33X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI33X0P7H7L A0 A1 A2 B0 B1 B2 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I B2:I Y:O VDD:B VSS:B
MMNM5 Y A2 net20 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM4 Y B2 net19 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM3 net20 A1 net21 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM2 net19 B1 net18 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM1 net21 A0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM0 net18 B0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMPM5 Y B1 net13 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM4 net13 A1 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM3 net13 A2 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM2 net13 A0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM1 Y B2 net13 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM0 Y B0 net13 VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI33X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI33X1H7L A0 A1 A2 B0 B1 B2 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I B2:I Y:O VDD:B VSS:B
MMNM5 Y A2 net20 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM4 Y B2 net19 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM3 net20 A1 net21 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM2 net19 B1 net18 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM1 net21 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM0 net18 B0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMPM5 Y B1 net13 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM4 net13 A1 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM3 net13 A2 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM2 net13 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM1 Y B2 net13 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM0 Y B0 net13 VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI33X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI33X1P4H7L A0 A1 A2 B0 B1 B2 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I B2:I Y:O VDD:B VSS:B
MMNM5 Y A2 net20 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM4 Y B2 net19 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM3 net20 A1 net21 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM2 net19 B1 net18 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM1 net21 A0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM0 net18 B0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMPM5 Y B1 net13 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM4 net13 A1 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM3 net13 A2 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM2 net13 A0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM1 Y B2 net13 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM0 Y B0 net13 VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI33X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI33X2H7L A0 A1 A2 B0 B1 B2 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I B2:I Y:O VDD:B VSS:B
MMPM4 net44 A1 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM5 Y B1 net44 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM3 net44 A2 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM0 Y B0 net44 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM1 Y B2 net44 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM2 net44 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMNM0 net42 B0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM1 net39 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM2 net41 B1 net42 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM3 net40 A1 net39 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM4 Y B2 net41 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM5 Y A2 net40 VSS nm1p2_lvt_lp W=300n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI33X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI33X3H7L A0 A1 A2 B0 B1 B2 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I B2:I Y:O VDD:B VSS:B
MMNM5 Y A2 net20 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM4 Y B2 net19 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM3 net20 A1 net21 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM2 net19 B1 net18 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM1 net21 A0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM0 net18 B0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMPM5 Y B1 net13 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM4 net13 A1 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM3 net13 A2 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM2 net13 A0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM1 Y B2 net13 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM0 Y B0 net13 VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    AOI33X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT AOI33X4H7L A0 A1 A2 B0 B1 B2 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I B2:I Y:O VDD:B VSS:B
MMNM5 Y A2 net20 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM4 Y B2 net19 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM3 net20 A1 net21 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM2 net19 B1 net18 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM1 net21 A0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM0 net18 B0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMPM5 Y B1 net13 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM4 net13 A1 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM3 net13 A2 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM2 net13 A0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM1 Y B2 net13 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM0 Y B0 net13 VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    BUFX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT BUFX0P5H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI1 net6 VDD VSS Y / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI0 A VDD VSS net6 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    BUFX0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT BUFX0P7H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI1 net6 VDD VSS Y / INV pl=6e-08 pw=2.22e-07 nl=6e-08 nw=1.74e-07
XXI0 A VDD VSS net6 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    BUFX10H7L
* View Name:    schematic
************************************************************************

.SUBCKT BUFX10H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI1 net6 VDD VSS Y / INV pl=6e-08 pw=19e-07 nl=6e-08 nw=15e-07
XXI0 A VDD VSS net6 / INV pl=6e-08 pw=7.6e-07 nl=6e-08 nw=6e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    BUFX12H7L
* View Name:    schematic
************************************************************************

.SUBCKT BUFX12H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI1 net6 VDD VSS Y / INV pl=6e-08 pw=2.28e-06 nl=6e-08 nw=1.8e-06
XXI0 A VDD VSS net6 / INV pl=6e-08 pw=9.3e-07 nl=6e-08 nw=7.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    BUFX16H7L
* View Name:    schematic
************************************************************************

.SUBCKT BUFX16H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI1 net6 VDD VSS Y / INV pl=6e-08 pw=3.04e-06 nl=6e-08 nw=2.4e-06
XXI0 A VDD VSS net6 / INV pl=6e-08 pw=1.14e-06 nl=6e-08 nw=9e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    BUFX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT BUFX1H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI1 net6 VDD VSS Y / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
XXI0 A VDD VSS net6 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    BUFX1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT BUFX1P4H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI1 net6 VDD VSS Y / INV pl=6e-08 pw=3.14e-07 nl=6e-08 nw=2.46e-07
XXI0 A VDD VSS net6 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    BUFX20H7L
* View Name:    schematic
************************************************************************

.SUBCKT BUFX20H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI1 net6 VDD VSS Y / INV pl=6e-08 pw=38e-07 nl=6e-08 nw=32e-07
XXI0 A VDD VSS net6 / INV pl=6e-08 pw=15.2e-07 nl=6e-08 nw=12e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    BUFX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT BUFX2H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI1 net6 VDD VSS Y / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
XXI0 A VDD VSS net6 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    BUFX2P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT BUFX2P5H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI1 net6 VDD VSS Y / INV pl=6e-08 pw=4.75e-07 nl=6e-08 nw=3.75e-07
XXI0 A VDD VSS net6 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    BUFX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT BUFX3H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI1 net6 VDD VSS Y / INV pl=6e-08 pw=5.7e-07 nl=6e-08 nw=4.5e-07
XXI0 A VDD VSS net6 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    BUFX3P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT BUFX3P5H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI1 net6 VDD VSS Y / INV pl=6e-08 pw=6.65e-07 nl=6e-08 nw=5.25e-07
XXI0 A VDD VSS net6 / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    BUFX4H7L
* View Name:    schematic
************************************************************************

.SUBCKT BUFX4H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI1 net6 VDD VSS Y / INV pl=6e-08 pw=7.6e-07 nl=6e-08 nw=6e-07
XXI0 A VDD VSS net6 / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    BUFX5H7L
* View Name:    schematic
************************************************************************

.SUBCKT BUFX5H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI1 net6 VDD VSS Y / INV pl=6e-08 pw=9.5e-07 nl=6e-08 nw=7.5e-07
XXI0 A VDD VSS net6 / INV pl=6e-08 pw=3.45e-07 nl=6e-08 nw=2.75e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    BUFX6H7L
* View Name:    schematic
************************************************************************

.SUBCKT BUFX6H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI0 A VDD VSS net4 / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
XXI1 net4 VDD VSS Y / INV pl=6e-08 pw=1.14e-06 nl=6e-08 nw=9e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    BUFX7H7L
* View Name:    schematic
************************************************************************

.SUBCKT BUFX7H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI1 net6 VDD VSS Y / INV pl=6e-08 pw=13.3e-07 nl=6e-08 nw=10.5e-07
XXI0 A VDD VSS net6 / INV pl=6e-08 pw=5e-07 nl=6e-08 nw=4e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    BUFX8H7L
* View Name:    schematic
************************************************************************

.SUBCKT BUFX8H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI0 A VDD VSS net4 / INV pl=6e-08 pw=6.2e-07 nl=6e-08 nw=5e-07
XXI1 net4 VDD VSS Y / INV pl=6e-08 pw=1.52e-06 nl=6e-08 nw=1.2e-06
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFNQX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFNQX1H7L CKN D Q VDD VSS
*.PININFO CKN:I D:I Q:O VDD:B VSS:B
XXI9 net73 net76 net71 VDD VSS net64 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI6 D net71 net76 VDD VSS net68 / TSINV pl=60n pw=200n nl=60n nw=160n
XXI15 net61 net71 net76 VDD VSS net64 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI14 net73 net76 net71 VDD VSS net68 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI4 CKN VDD VSS net76 / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI7 net68 VDD VSS net73 / INV pl=60n pw=190n nl=60n nw=150n
XXI13 net76 VDD VSS net71 / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI12 net64 VDD VSS Q / INV pl=60n pw=270n nl=60n nw=210n
XXI10 net64 VDD VSS net61 / INV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFNQX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFNQX2H7L CKN D Q VDD VSS
*.PININFO CKN:I D:I Q:O VDD:B VSS:B
XXI9 net73 net76 net71 VDD VSS net64 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI6 D net71 net76 VDD VSS net68 / TSINV pl=60n pw=210n nl=60n nw=170n
XXI15 net61 net71 net76 VDD VSS net64 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI14 net73 net76 net71 VDD VSS net68 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI4 CKN VDD VSS net76 / INV pl=60n pw=210n nl=60n nw=170n
XXI7 net68 VDD VSS net73 / INV pl=60n pw=200n nl=60n nw=160n
XXI13 net76 VDD VSS net71 / INV pl=60n pw=210n nl=60n nw=170n
XXI12 net64 VDD VSS Q / INV pl=60n pw=380n nl=60n nw=300n
XXI10 net64 VDD VSS net61 / INV pl=60n pw=210n nl=60n nw=170n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFNQX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFNQX3H7L CKN D Q VDD VSS
*.PININFO CKN:I D:I Q:O VDD:B VSS:B
XXI9 net73 net76 net71 VDD VSS net64 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI6 D net71 net76 VDD VSS net68 / TSINV pl=60n pw=220n nl=60n nw=175n
XXI15 net61 net71 net76 VDD VSS net64 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI14 net73 net76 net71 VDD VSS net68 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI4 CKN VDD VSS net76 / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI7 net68 VDD VSS net73 / INV pl=60n pw=205n nl=60n nw=165n
XXI13 net76 VDD VSS net71 / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI12 net64 VDD VSS Q / INV pl=60n pw=570n nl=60n nw=450n
XXI10 net64 VDD VSS net61 / INV pl=60n pw=230n nl=60n nw=185n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFNRX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFNRX0P5H7L CKN D Q QN RN VDD VSS
*.PININFO CKN:I D:I RN:I Q:O QN:O VDD:B VSS:B
MMN1 net085 CKB net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0124 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net085 R VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN4 net46 net33 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMP4 net54 R VDD VDD pm1p2_lvt_lp W=280n L=60n m=1
MMP2 net67 net0124 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net085 CKP net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=280n L=60n m=1
XXI29 net46 CKP CKB VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XI3 D CKB CKP VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2.4E-07
XI6 net085 VDD VSS QN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI2 RN VDD VSS R / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI5 net0124 VDD VSS Q / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI1 CKP VDD VSS CKB / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI4 net085 VDD VSS net0124 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI0 CKN VDD VSS CKP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI9 CKP CKB net46 net085 VDD VSS / TG pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFNRX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFNRX1H7L CKN D Q QN RN VDD VSS
*.PININFO CKN:I D:I RN:I Q:O QN:O VDD:B VSS:B
MMN1 net085 CKB net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0124 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net085 R VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN4 net46 net33 VSS VSS nm1p2_lvt_lp W=220n L=60n m=1
MMP4 net54 R VDD VDD pm1p2_lvt_lp W=300n L=60n m=1
MMP2 net67 net0124 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net085 CKP net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=300n L=60n m=1
XXI29 net46 CKP CKB VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XI3 D CKB CKP VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2.4E-07
XI7 net085 VDD VSS QN / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI2 RN VDD VSS R / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI5 net0124 VDD VSS Q / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI1 CKP VDD VSS CKB / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI4 net085 VDD VSS net0124 / INV pl=6E-08 pw=3E-07 nl=6E-08 nw=2.2E-07
XI0 CKN VDD VSS CKP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI9 CKP CKB net46 net085 VDD VSS / TG pl=6E-08 pw=3E-07 nl=6E-08 nw=2.2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFNRX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFNRX2H7L CKN D Q QN RN VDD VSS
*.PININFO CKN:I D:I RN:I Q:O QN:O VDD:B VSS:B
MMN1 net085 CKB net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0124 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net085 R VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN4 net46 net33 VSS VSS nm1p2_lvt_lp W=240n L=60n m=1
MMP4 net54 R VDD VDD pm1p2_lvt_lp W=340n L=60n m=1
MMP2 net67 net0124 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net085 CKP net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=340n L=60n m=1
XXI29 net46 CKP CKB VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XI3 D CKB CKP VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2.4E-07
XI10 net085 VDD VSS QN / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI7 CKP VDD VSS CKB / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI5 net0124 VDD VSS Q / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI8 RN VDD VSS R / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI9 net085 VDD VSS net0124 / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI0 CKN VDD VSS CKP / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI9 CKP CKB net46 net085 VDD VSS / TG pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFNRX4H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFNRX4H7L CKN D Q QN RN VDD VSS
*.PININFO CKN:I D:I RN:I Q:O QN:O VDD:B VSS:B
MMN1 net085 CKB net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0124 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net085 R VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN4 net46 net33 VSS VSS nm1p2_lvt_lp W=260n L=60n m=1
MMP4 net54 R VDD VDD pm1p2_lvt_lp W=360n L=60n m=1
MMP2 net67 net0124 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net085 CKP net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=360n L=60n m=1
XXI29 net46 CKP CKB VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XI3 D CKB CKP VDD VSS net33 / TSINV pl=6E-08 pw=3.2E-07 nl=6E-08 nw=2.6E-07
XI11 net085 VDD VSS QN / INV pl=6E-08 pw=8E-07 nl=6E-08 nw=5.6E-07
XI7 CKP VDD VSS CKB / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI5 net0124 VDD VSS Q / INV pl=6E-08 pw=8E-07 nl=6E-08 nw=5.6E-07
XI8 RN VDD VSS R / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI9 net085 VDD VSS net0124 / INV pl=6E-08 pw=3.6E-07 nl=6E-08 nw=2.6E-07
XI0 CKN VDD VSS CKP / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI9 CKP CKB net46 net085 VDD VSS / TG pl=6E-08 pw=3.35E-07 nl=6E-08 nw=2.6E-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFNSRQX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFNSRQX1H7L CKN D Q RN SN VDD VSS
*.PININFO CKN:I D:I RN:I SN:I Q:O VDD:B VSS:B
XI3 net0144 VDD VSS Q / INV pl=6E-08 pw=2.7E-07 nl=6E-08 nw=2.1E-07
XI2 net094 VDD VSS net0144 / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XI1 RN VDD VSS R / INV pl=6E-08 pw=1.7E-07 nl=6E-08 nw=1.5E-07
XI0 CKP VDD VSS CKB / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI4 CKN VDD VSS CKP / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI30 D CKB CKP VDD VSS net33 / TSINV pl=6E-08 pw=2E-07 nl=6E-08 nw=1.6E-07
XXI29 net46 CKP CKB VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
MMN6 net094 R net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 net062 VSS nm1p2_lvt_lp W=170n L=60n m=1
MMN1 net094 CKB net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0144 net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net062 SN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
XXI9 CKP CKB net46 net094 VDD VSS / TG pl=6E-08 pw=1.5E-07 nl=6E-08 nw=1.5E-07
MMP5 net54 R VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP2 net67 net0144 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=210n L=60n m=1
MMP4 net094 SN VDD VDD pm1p2_lvt_lp W=170n L=60n m=1
MMP1 net094 CKP net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFNSRQX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFNSRQX2H7L CKN D Q RN SN VDD VSS
*.PININFO CKN:I D:I RN:I SN:I Q:O VDD:B VSS:B
XI3 net0144 VDD VSS Q / INV pl=6E-08 pw=3.8E-07 nl=6E-08 nw=3E-07
XI2 net094 VDD VSS net0144 / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XI1 RN VDD VSS R / INV pl=6E-08 pw=1.5E-07 nl=6E-08 nw=1.5E-07
XI0 CKP VDD VSS CKB / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI4 CKN VDD VSS CKP / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI30 D CKB CKP VDD VSS net33 / TSINV pl=6E-08 pw=2E-07 nl=6E-08 nw=1.6E-07
XXI29 net46 CKP CKB VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
MMN6 net094 R net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 net062 VSS nm1p2_lvt_lp W=170n L=60n m=1
MMN1 net094 CKB net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0144 net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net062 SN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
XXI9 CKP CKB net46 net094 VDD VSS / TG pl=6E-08 pw=1.9E-07 nl=6E-08 nw=1.5E-07
MMP5 net54 R VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP2 net67 net0144 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=210n L=60n m=1
MMP4 net094 SN VDD VDD pm1p2_lvt_lp W=180n L=60n m=1
MMP1 net094 CKP net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFNSRX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFNSRX0P5H7L CKN D Q QN RN SN VDD VSS
*.PININFO CKN:I D:I RN:I SN:I Q:O QN:O VDD:B VSS:B
XI3 net0144 VDD VSS Q / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI2 net094 VDD VSS net0144 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI1 RN VDD VSS R / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI4 net094 VDD VSS QN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI0 CKP VDD VSS CKB / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI4 CKN VDD VSS CKP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI30 D CKB CKP VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI29 net46 CKP CKB VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
MMN4 net46 net33 net062 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN1 net094 CKB net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN6 net094 R net062 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN2 net36 net0144 net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net062 SN VSS VSS nm1p2_lvt_lp W=240n L=60n m=1
XXI9 CKP CKB net46 net094 VDD VSS / TG pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
MMP5 net54 R VDD VDD pm1p2_lvt_lp W=280n L=60n m=1
MMP2 net67 net0144 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP4 net094 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=280n L=60n m=1
MMP1 net094 CKP net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFNSRX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFNSRX1H7L CKN D Q QN RN SN VDD VSS
*.PININFO CKN:I D:I RN:I SN:I Q:O QN:O VDD:B VSS:B
XI3 net0144 VDD VSS Q / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI2 net094 VDD VSS net0144 / INV pl=6E-08 pw=3E-07 nl=6E-08 nw=2.2E-07
XI1 RN VDD VSS R / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI5 net094 VDD VSS QN / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI0 CKP VDD VSS CKB / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI4 CKN VDD VSS CKP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI30 D CKB CKP VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI29 net46 CKP CKB VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
MMN6 net094 R net062 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN4 net46 net33 net062 VSS nm1p2_lvt_lp W=215n L=60n m=1
MMN1 net094 CKB net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0144 net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net062 SN VSS VSS nm1p2_lvt_lp W=240n L=60n m=1
XXI9 CKP CKB net46 net094 VDD VSS / TG pl=6E-08 pw=3E-07 nl=6E-08 nw=2.2E-07
MMP5 net54 R VDD VDD pm1p2_lvt_lp W=300n L=60n m=1
MMP2 net67 net0144 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=300n L=60n m=1
MMP4 net094 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP1 net094 CKP net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFNSRX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFNSRX2H7L CKN D Q QN RN SN VDD VSS
*.PININFO CKN:I D:I RN:I SN:I Q:O QN:O VDD:B VSS:B
XI3 net0144 VDD VSS Q / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI8 net094 VDD VSS net0144 / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI6 RN VDD VSS R / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI7 net094 VDD VSS QN / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI5 CKP VDD VSS CKB / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI4 CKN VDD VSS CKP / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI30 D CKB CKP VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI29 net46 CKP CKB VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
MMN6 net094 R net062 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN4 net46 net33 net062 VSS nm1p2_lvt_lp W=240n L=60n m=1
MMN1 net094 CKB net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0144 net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net062 SN VSS VSS nm1p2_lvt_lp W=260n L=60n m=1
XXI9 CKP CKB net46 net094 VDD VSS / TG pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
MMP5 net54 R VDD VDD pm1p2_lvt_lp W=340n L=60n m=1
MMP2 net67 net0144 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=340n L=60n m=1
MMP4 net094 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP1 net094 CKP net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFNSX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFNSX0P5H7L CKN D Q QN SN VDD VSS
*.PININFO CKN:I D:I SN:I Q:O QN:O VDD:B VSS:B
MMN6 net056 SN VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMN1 net082 CKB net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net048 net056 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 net056 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMP0 net082 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP2 net67 net048 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net082 CKP net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 VDD VDD pm1p2_lvt_lp W=280n L=60n m=1
XI0 D CKB CKP VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI1 net46 CKP CKB VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08 nw=1.5E-07
XI5 net082 VDD VSS net048 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI4 net048 VDD VSS Q / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI2 CKP VDD VSS CKB / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI3 net082 VDD VSS QN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI4 CKN VDD VSS CKP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI9 CKP CKB net46 net082 VDD VSS / TG pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFNSX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFNSX1H7L CKN D Q QN SN VDD VSS
*.PININFO CKN:I D:I SN:I Q:O QN:O VDD:B VSS:B
MMN6 net056 SN VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMN1 net082 CKB net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net048 net056 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 net056 VSS nm1p2_lvt_lp W=220n L=60n m=1
MMP0 net082 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP2 net67 net048 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net082 CKP net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 VDD VDD pm1p2_lvt_lp W=300n L=60n m=1
XI0 D CKB CKP VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI1 net46 CKP CKB VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08 nw=1.5E-07
XI5 net082 VDD VSS net048 / INV pl=6E-08 pw=3E-07 nl=6E-08 nw=2.2E-07
XI4 net048 VDD VSS Q / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI2 CKP VDD VSS CKB / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI6 net082 VDD VSS QN / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI4 CKN VDD VSS CKP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI9 CKP CKB net46 net082 VDD VSS / TG pl=6E-08 pw=3E-07 nl=6E-08 nw=2.2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFNSX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFNSX2H7L CKN D Q QN SN VDD VSS
*.PININFO CKN:I D:I SN:I Q:O QN:O VDD:B VSS:B
MMN6 net056 SN VSS VSS nm1p2_lvt_lp W=240n L=60n m=1
MMN1 net082 CKB net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net048 net056 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 net056 VSS nm1p2_lvt_lp W=240n L=60n m=1
MMP0 net082 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP2 net67 net048 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net082 CKP net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 VDD VDD pm1p2_lvt_lp W=340n L=60n m=1
XI0 D CKB CKP VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI1 net46 CKP CKB VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08 nw=1.5E-07
XI7 net082 VDD VSS net048 / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI8 net048 VDD VSS Q / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI6 CKP VDD VSS CKB / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI3 net082 VDD VSS QN / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XXI4 CKN VDD VSS CKP / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI9 CKP CKB net46 net082 VDD VSS / TG pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFNX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFNX0P5H7L CKN D Q QN VDD VSS
*.PININFO CKN:I D:I Q:O QN:O VDD:B VSS:B
XI3 net61 CKB CKP VDD VSS net64 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08 nw=1.5E-07
XXI29 net73 CKP CKB VDD VSS net68 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI30 D CKB CKP VDD VSS net68 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI4 net73 CKP CKB VDD VSS net64 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI7 net64 VDD VSS Q / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI5 net64 VDD VSS net61 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI6 net61 VDD VSS QN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI1 CKP VDD VSS CKB / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI2 net68 VDD VSS net73 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI0 CKN VDD VSS CKP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFNX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFNX1H7L CKN D Q QN VDD VSS
*.PININFO CKN:I D:I Q:O QN:O VDD:B VSS:B
XI3 net61 CKB CKP VDD VSS net64 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08 nw=1.5E-07
XXI29 net73 CKP CKB VDD VSS net68 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI30 D CKB CKP VDD VSS net68 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI4 net73 CKP CKB VDD VSS net64 / TSINV pl=6E-08 pw=3E-07 nl=6E-08 nw=2.2E-07
XI8 net64 VDD VSS Q / INV pl=6E-08 pw=3E-07 nl=6E-08 nw=2.4E-07
XI5 net64 VDD VSS net61 / INV pl=6E-08 pw=3E-07 nl=6E-08 nw=2.2E-07
XI6 net61 VDD VSS QN / INV pl=6E-08 pw=3E-07 nl=6E-08 nw=2.4E-07
XI1 CKP VDD VSS CKB / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI2 net68 VDD VSS net73 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI0 CKN VDD VSS CKP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFNX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFNX2H7L CKN D Q QN VDD VSS
*.PININFO CKN:I D:I Q:O QN:O VDD:B VSS:B
XI9 D CKB CKP VDD VSS net68 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI3 net61 CKB CKP VDD VSS net64 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08 nw=1.5E-07
XXI29 net73 CKP CKB VDD VSS net68 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XI4 net73 CKP CKB VDD VSS net64 / TSINV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI12 net64 VDD VSS Q / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI11 net64 VDD VSS net61 / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI6 net61 VDD VSS QN / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI8 CKP VDD VSS CKB / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI10 net68 VDD VSS net73 / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI0 CKN VDD VSS CKP / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFNX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFNX3H7L CKN D Q QN VDD VSS
*.PININFO CKN:I D:I Q:O QN:O VDD:B VSS:B
XI4 net73 CKP CKB VDD VSS net64 / TSINV pl=60n pw=360n nl=60n nw=260n
XXI29 net73 CKP CKB VDD VSS net68 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XI3 net61 CKB CKP VDD VSS net64 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08 nw=1.5E-07
XI9 D CKB CKP VDD VSS net68 / TSINV pl=60n pw=340n nl=60n nw=240n
XI0 CKN VDD VSS CKP / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI10 net68 VDD VSS net73 / INV pl=60n pw=360n nl=60n nw=260n
XI8 CKP VDD VSS CKB / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI6 net61 VDD VSS QN / INV pl=60n pw=600n nl=60n nw=420n
XI11 net64 VDD VSS net61 / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI12 net64 VDD VSS Q / INV pl=60n pw=600n nl=60n nw=420n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFQX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFQX0P5H7L CK D Q VDD VSS
*.PININFO CK:I D:I Q:O VDD:B VSS:B
XXI14 net46 net24 net32 VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI6 D net32 net24 VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI9 net46 net24 net32 VDD VSS net25 / TSINV pl=6E-08 pw=3.2E-07 nl=6E-08
+ nw=2.3E-07
XXI15 net9 net32 net24 VDD VSS net25 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI7 net33 VDD VSS net46 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI13 net32 VDD VSS net24 / INV pl=6E-08 pw=3.1E-07 nl=6E-08 nw=2.2E-07
XXI12 net25 VDD VSS Q / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI10 net25 VDD VSS net9 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI4 CK VDD VSS net32 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFQX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFQX1H7L CK D Q VDD VSS
*.PININFO CK:I D:I Q:O VDD:B VSS:B
XXI14 net46 net24 net32 VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI6 D net32 net24 VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI9 net46 net24 net32 VDD VSS net25 / TSINV pl=6E-08 pw=3.2E-07 nl=6E-08
+ nw=2.3E-07
XXI15 net9 net32 net24 VDD VSS net25 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI7 net33 VDD VSS net46 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI13 net32 VDD VSS net24 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI12 net25 VDD VSS Q / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI10 net25 VDD VSS net9 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI4 CK VDD VSS net32 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFQX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFQX2H7L CK D Q VDD VSS
*.PININFO CK:I D:I Q:O VDD:B VSS:B
XXI14 net46 net24 net32 VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI6 D net32 net24 VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI9 net46 net24 net32 VDD VSS net25 / TSINV pl=6E-08 pw=3.4E-07 nl=6E-08
+ nw=2.4E-07
XXI15 net9 net32 net24 VDD VSS net25 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI7 net33 VDD VSS net46 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI13 net32 VDD VSS net24 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI12 net25 VDD VSS Q / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XXI10 net25 VDD VSS net9 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI4 CK VDD VSS net32 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFQX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFQX3H7L CK D Q VDD VSS
*.PININFO CK:I D:I Q:O VDD:B VSS:B
XXI14 net46 net24 net32 VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI6 D net32 net24 VDD VSS net33 / TSINV pl=6E-08 pw=3.1E-07 nl=6E-08
+ nw=2.2E-07
XXI9 net46 net24 net32 VDD VSS net25 / TSINV pl=6E-08 pw=3.1E-07 nl=6E-08
+ nw=2.2E-07
XXI15 net9 net32 net24 VDD VSS net25 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI7 net33 VDD VSS net46 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI13 net32 VDD VSS net24 / INV pl=6E-08 pw=3.1E-07 nl=6E-08 nw=2.2E-07
XXI12 net25 VDD VSS Q / INV pl=6E-08 pw=6E-07 nl=6E-08 nw=4.2E-07
XXI10 net25 VDD VSS net9 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI4 CK VDD VSS net32 / INV pl=6E-08 pw=3.1E-07 nl=6E-08 nw=2.2E-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net15 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 net15 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP2 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFRQNX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFRQNX1H7L CK D QN RN VDD VSS
*.PININFO CK:I D:I RN:I QN:O VDD:B VSS:B
MMM19 net40 cn net33 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM18 net33 net25 net61 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM28 net61 RN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM22 net40 c net117 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMM21 net117 net25 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMM27 net117 RN VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
XXI6 CK VDD VSS cn / INV pl=60n pw=210n nl=60n nw=170n
XXI5 cn VDD VSS c / INV pl=60n pw=210n nl=60n nw=170n
XI2 D VDD VSS net53 / INV pl=60n pw=190n nl=60n nw=150n
XI6 net25 VDD VSS QN / INV pl=60n pw=270n nl=60n nw=210n
XI4 net40 VDD VSS net25 / INV pl=60n pw=190n nl=60n nw=150n
XI3 net51 c cn VDD VSS net13 / TSINV pl=60n pw=150n nl=60n nw=150n
XI7 net53 cn c VDD VSS net13 / TSINV pl=60n pw=200n nl=60n nw=240n
XI0 RN net13 VDD VSS net51 / NAND2 pl=60n pw=210n nl=60n nw=170n
XI5 c cn net51 net40 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net15 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 net15 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP2 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFRQNX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFRQNX2H7L CK D QN RN VDD VSS
*.PININFO CK:I D:I RN:I QN:O VDD:B VSS:B
MNM2 net72 RN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net71 net25 net72 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net40 cn net71 VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM1 net70 net25 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM2 net70 RN VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM0 net40 c net70 VDD pm1p2_lvt_lp W=150n L=60n m=1
XXI5 cn VDD VSS c / INV pl=60n pw=210n nl=60n nw=170n
XXI6 CK VDD VSS cn / INV pl=60n pw=210n nl=60n nw=170n
XI2 D VDD VSS net53 / INV pl=60n pw=190n nl=60n nw=150n
XI4 net40 VDD VSS net25 / INV pl=60n pw=210n nl=60n nw=170n
XI6 net25 VDD VSS QN / INV pl=60n pw=380n nl=60n nw=300n
XI3 net51 c cn VDD VSS net13 / TSINV pl=60n pw=150n nl=60n nw=150n
XI7 net53 cn c VDD VSS net13 / TSINV pl=60n pw=200n nl=60n nw=240n
XI0 RN net13 VDD VSS net51 / NAND2 pl=60n pw=210n nl=60n nw=170n
XI5 c cn net51 net40 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net15 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 net15 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP2 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFRQX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFRQX0P5H7L CK D Q RN VDD VSS
*.PININFO CK:I D:I RN:I Q:O VDD:B VSS:B
MMN1 net43 net41 net40 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net40 RN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 net46 net71 net43 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP2 net46 RN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP1 net55 net41 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP0 net46 net63 net55 VDD pm1p2_lvt_lp W=150n L=60n m=1
XXI21 net66 net63 net71 VDD VSS net61 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI6 net77 net71 net63 VDD VSS net61 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08
+ nw=2.4E-07
XXI20 RN net61 VDD VSS net66 / NAND2 pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2.4E-07
XXI19 net46 VDD VSS net41 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI23 D VDD VSS net77 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI13 net71 VDD VSS net63 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI26 net46 VDD VSS Q / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI4 CK VDD VSS net71 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI22 net63 net71 net66 net46 VDD VSS / TG pl=6E-08 pw=2.8E-07 nl=6E-08
+ nw=2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net15 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 net15 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP2 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFRQX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFRQX1H7L CK D Q RN VDD VSS
*.PININFO CK:I D:I RN:I Q:O VDD:B VSS:B
MMN0 net55 net71 net43 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net40 RN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 net43 net41 net40 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP2 net55 RN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP0 net55 net63 net049 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net049 net41 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
XXI21 net66 net63 net71 VDD VSS net61 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI6 net77 net71 net63 VDD VSS net61 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08
+ nw=2.4E-07
XXI20 RN net61 VDD VSS net66 / NAND2 pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2.4E-07
XXI23 D VDD VSS net77 / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI19 net55 VDD VSS net41 / INV pl=6E-08 pw=3E-07 nl=6E-08 nw=2.2E-07
XXI13 net71 VDD VSS net63 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI26 net55 VDD VSS Q / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI4 CK VDD VSS net71 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI22 net63 net71 net66 net55 VDD VSS / TG pl=6E-08 pw=3E-07 nl=6E-08
+ nw=2.2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net15 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 net15 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP2 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFRQX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFRQX2H7L CK D Q RN VDD VSS
*.PININFO CK:I D:I RN:I Q:O VDD:B VSS:B
MMN2 net40 RN VSS VSS nm1p2_lvt_lp W=260n L=60n m=1
MMN0 net46 net71 net43 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 net43 net41 net40 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP2 net46 RN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP0 net46 net63 net49 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net49 net41 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
XXI21 net66 net63 net71 VDD VSS net61 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI6 net77 net71 net63 VDD VSS net61 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08
+ nw=2.4E-07
XXI20 RN net61 VDD VSS net66 / NAND2 pl=6E-08 pw=2E-07 nl=6E-08 nw=2.4E-07
XXI23 D VDD VSS net77 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2.4E-07
XXI4 CK VDD VSS net71 / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI19 net46 VDD VSS net41 / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI26 net46 VDD VSS Q / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XXI13 net71 VDD VSS net63 / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI22 net63 net71 net66 net46 VDD VSS / TG pl=6E-08 pw=3.4E-07 nl=6E-08
+ nw=2.4E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFRX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFRX0P5H7L CK D Q QN RN VDD VSS
*.PININFO CK:I D:I RN:I Q:O QN:O VDD:B VSS:B
MNM0 net36 net0122 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 net042 CKN net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net042 R VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN4 net46 net33 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMP4 net54 R VDD VDD pm1p2_lvt_lp W=280n L=60n m=1
MMP1 net042 CKP net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=280n L=60n m=1
MPM0 net67 net0122 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
XXI29 net46 CKP CKN VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI30 D CKN CKP VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2.4E-07
XI3 net042 VDD VSS QN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI1 RN VDD VSS R / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI4 net0122 VDD VSS Q / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI0 CKN VDD VSS CKP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI2 net042 VDD VSS net0122 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI4 CK VDD VSS CKN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI9 CKP CKN net46 net042 VDD VSS / TG pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFRX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFRX1H7L CK D Q QN RN VDD VSS
*.PININFO CK:I D:I RN:I Q:O QN:O VDD:B VSS:B
MNM0 net36 net0122 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 net042 CKN net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net042 R VSS VSS nm1p2_lvt_lp W=220n L=60n m=1
MMN4 net46 net33 VSS VSS nm1p2_lvt_lp W=220n L=60n m=1
MMP4 net54 R VDD VDD pm1p2_lvt_lp W=300n L=60n m=1
MMP1 net042 CKP net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=300n L=60n m=1
MPM0 net67 net0122 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
XXI29 net46 CKP CKN VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI30 D CKN CKP VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2.4E-07
XI3 net042 VDD VSS QN / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI1 RN VDD VSS R / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI5 net0122 VDD VSS Q / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI0 CKN VDD VSS CKP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI2 net042 VDD VSS net0122 / INV pl=6E-08 pw=3E-07 nl=6E-08 nw=2.2E-07
XXI4 CK VDD VSS CKN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI9 CKP CKN net46 net042 VDD VSS / TG pl=6E-08 pw=3E-07 nl=6E-08 nw=2.2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFRX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFRX2H7L CK D Q QN RN VDD VSS
*.PININFO CK:I D:I RN:I Q:O QN:O VDD:B VSS:B
MNM0 net36 net0122 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 net042 CKN net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net042 R VSS VSS nm1p2_lvt_lp W=240n L=60n m=1
MMN4 net46 net33 VSS VSS nm1p2_lvt_lp W=240n L=60n m=1
MMP4 net54 R VDD VDD pm1p2_lvt_lp W=340n L=60n m=1
MMP1 net042 CKP net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=340n L=60n m=1
MPM0 net67 net0122 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
XXI30 D CKN CKP VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2.4E-07
XXI29 net46 CKP CKN VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XI8 net042 VDD VSS net0122 / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI6 CKN VDD VSS CKP / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI9 net0122 VDD VSS Q / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI7 RN VDD VSS R / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI3 net042 VDD VSS QN / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI5 CK VDD VSS CKN / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI9 CKP CKN net46 net042 VDD VSS / TG pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFRX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFRX3H7L CK D Q QN RN VDD VSS
*.PININFO CK:I D:I RN:I Q:O QN:O VDD:B VSS:B
MNM0 net17 net0122 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 net042 CKN net17 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net042 R VSS VSS nm1p2_lvt_lp W=260n L=60n m=1
MMN4 net46 net33 VSS VSS nm1p2_lvt_lp W=260n L=60n m=1
MMP4 net92 R VDD VDD pm1p2_lvt_lp W=360n L=60n m=1
MMP1 net042 CKP net25 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net92 VDD pm1p2_lvt_lp W=360n L=60n m=1
MPM0 net25 net0122 net92 VDD pm1p2_lvt_lp W=150n L=60n m=1
XXI29 net46 CKP CKN VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI30 D CKN CKP VDD VSS net33 / TSINV pl=60n pw=320n nl=60n nw=260n
XI5 CK VDD VSS CKN / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI3 net042 VDD VSS QN / INV pl=60n pw=600n nl=60n nw=420n
XI7 RN VDD VSS R / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI9 net0122 VDD VSS Q / INV pl=60n pw=600n nl=60n nw=420n
XI6 CKN VDD VSS CKP / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI8 net042 VDD VSS net0122 / INV pl=60n pw=360n nl=60n nw=260n
XXI9 CKP CKN net46 net042 VDD VSS / TG pl=60n pw=360n nl=60n nw=260n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFSQNX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFSQNX1H7L CK D QN SN VDD VSS
*.PININFO CK:I D:I SN:I QN:O VDD:B VSS:B
MMN1 net0161 net32 net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net048 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net0161 net086 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net087 net33 VSS VSS nm1p2_lvt_lp W=190n L=60n m=1
MMP4 net54 net086 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP2 net058 net048 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net0161 net24 net058 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net087 net33 net54 VDD pm1p2_lvt_lp W=200n L=60n m=1
XXI29 net087 net24 net32 VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI30 net080 net32 net24 VDD VSS net33 / TSINV pl=6E-08 pw=2E-07 nl=6E-08
+ nw=2E-07
XXI37 D VDD VSS net080 / INV pl=6E-08 pw=2.7E-07 nl=6E-08 nw=2.1E-07
XXI12 net048 VDD VSS QN / INV pl=6E-08 pw=2.7E-07 nl=6E-08 nw=2.1E-07
XXI31 SN VDD VSS net086 / INV pl=6E-08 pw=1.5E-07 nl=6E-08 nw=1.5E-07
XXI13 net32 VDD VSS net24 / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI10 net0161 VDD VSS net048 / INV pl=6E-08 pw=1.9E-07 nl=6E-08 nw=1.5E-07
XXI4 CK VDD VSS net32 / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI9 net24 net32 net087 net0161 VDD VSS / TG pl=6E-08 pw=1.9E-07 nl=6E-08
+ nw=1.5E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFSQNX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFSQNX2H7L CK D QN SN VDD VSS
*.PININFO CK:I D:I SN:I QN:O VDD:B VSS:B
MMN1 net0161 net32 net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net048 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net0161 net086 VSS VSS nm1p2_lvt_lp W=190n L=60n m=1
MMN4 net087 net33 VSS VSS nm1p2_lvt_lp W=190n L=60n m=1
MMP4 net54 net086 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP2 net059 net048 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net0161 net24 net059 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net087 net33 net54 VDD pm1p2_lvt_lp W=200n L=60n m=1
XXI29 net087 net24 net32 VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI30 net082 net32 net24 VDD VSS net33 / TSINV pl=6E-08 pw=2.1E-07 nl=6E-08
+ nw=2.1E-07
XXI38 D VDD VSS net082 / INV pl=6E-08 pw=3.8E-07 nl=6E-08 nw=3E-07
XXI12 net048 VDD VSS QN / INV pl=6E-08 pw=3.8E-07 nl=6E-08 nw=3E-07
XXI31 SN VDD VSS net086 / INV pl=6E-08 pw=1.5E-07 nl=6E-08 nw=1.5E-07
XXI13 net32 VDD VSS net24 / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI10 net0161 VDD VSS net048 / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI4 CK VDD VSS net32 / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI9 net24 net32 net087 net0161 VDD VSS / TG pl=6E-08 pw=1.9E-07 nl=6E-08
+ nw=1.5E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFSQX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFSQX1H7L CK D Q SN VDD VSS
*.PININFO CK:I D:I SN:I Q:O VDD:B VSS:B
MMN1 net0161 net32 net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net048 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net0161 net086 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net087 net33 VSS VSS nm1p2_lvt_lp W=190n L=60n m=1
MMP4 net54 net086 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP2 net058 net048 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net0161 net24 net058 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net087 net33 net54 VDD pm1p2_lvt_lp W=200n L=60n m=1
XXI29 net087 net24 net32 VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI30 net080 net32 net24 VDD VSS net33 / TSINV pl=6E-08 pw=2E-07 nl=6E-08
+ nw=2E-07
XXI37 D VDD VSS net080 / INV pl=6E-08 pw=2.7E-07 nl=6E-08 nw=2.1E-07
XXI12 net0161 VDD VSS Q / INV pl=6E-08 pw=2.7E-07 nl=6E-08 nw=2.1E-07
XXI31 SN VDD VSS net086 / INV pl=6E-08 pw=1.5E-07 nl=6E-08 nw=1.5E-07
XXI13 net32 VDD VSS net24 / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI10 net0161 VDD VSS net048 / INV pl=6E-08 pw=1.9E-07 nl=6E-08 nw=1.5E-07
XXI4 CK VDD VSS net32 / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI9 net24 net32 net087 net0161 VDD VSS / TG pl=6E-08 pw=1.9E-07 nl=6E-08
+ nw=1.5E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFSQX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFSQX2H7L CK D Q SN VDD VSS
*.PININFO CK:I D:I SN:I Q:O VDD:B VSS:B
MMN1 net0161 net32 net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net048 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net0161 net086 VSS VSS nm1p2_lvt_lp W=190n L=60n m=1
MMN4 net087 net33 VSS VSS nm1p2_lvt_lp W=190n L=60n m=1
MMP4 net54 net086 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP2 net059 net048 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net0161 net24 net059 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net087 net33 net54 VDD pm1p2_lvt_lp W=200n L=60n m=1
XXI29 net087 net24 net32 VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI30 net082 net32 net24 VDD VSS net33 / TSINV pl=6E-08 pw=2.1E-07 nl=6E-08
+ nw=2.1E-07
XXI38 D VDD VSS net082 / INV pl=6E-08 pw=3.8E-07 nl=6E-08 nw=3E-07
XXI12 net0161 VDD VSS Q / INV pl=6E-08 pw=3.8E-07 nl=6E-08 nw=3E-07
XXI31 SN VDD VSS net086 / INV pl=6E-08 pw=1.5E-07 nl=6E-08 nw=1.5E-07
XXI13 net32 VDD VSS net24 / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI10 net0161 VDD VSS net048 / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI4 CK VDD VSS net32 / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI9 net24 net32 net087 net0161 VDD VSS / TG pl=6E-08 pw=1.9E-07 nl=6E-08
+ nw=1.5E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFSRQX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFSRQX1H7L CK D Q RN SN VDD VSS
*.PININFO CK:I D:I RN:I SN:I Q:O VDD:B VSS:B
MMN5 net062 SN VSS VSS nm1p2_lvt_lp W=190n L=60n m=1
MMN1 net094 net0108 net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0144 net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN6 net094 net096 net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 net062 VSS nm1p2_lvt_lp W=190n L=60n m=1
MMP4 net094 SN VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP5 net54 net096 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP2 net67 net0144 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net094 net24 net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=200n L=60n m=1
XXI29 net46 net24 net0108 VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI30 D net0108 net24 VDD VSS net33 / TSINV pl=6E-08 pw=2E-07 nl=6E-08
+ nw=2.1E-07
XXI32 RN VDD VSS net096 / INV pl=6E-08 pw=1.5E-07 nl=6E-08 nw=1.5E-07
XXI5 net0144 VDD VSS Q / INV pl=6E-08 pw=2.7E-07 nl=6E-08 nw=2.1E-07
XXI13 net0108 VDD VSS net24 / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI10 net094 VDD VSS net0144 / INV pl=6E-08 pw=1.9E-07 nl=6E-08 nw=1.5E-07
XXI4 CK VDD VSS net0108 / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI9 net24 net0108 net46 net094 VDD VSS / TG pl=6E-08 pw=1.9E-07 nl=6E-08
+ nw=1.5E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFSRQX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFSRQX2H7L CK D Q RN SN VDD VSS
*.PININFO CK:I D:I RN:I SN:I Q:O VDD:B VSS:B
MMN5 net062 SN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 net0122 net0106 net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0143 net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP0 net0122 net096 net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 net062 VSS nm1p2_lvt_lp W=190n L=60n m=1
MMP4 net0122 SN VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP5 net54 net096 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP2 net67 net0143 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net0122 net24 net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=200n L=60n m=1
XXI29 net46 net24 net0106 VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI30 D net0106 net24 VDD VSS net33 / TSINV pl=6E-08 pw=2E-07 nl=6E-08
+ nw=2.1E-07
XXI32 RN VDD VSS net096 / INV pl=6E-08 pw=1.5E-07 nl=6E-08 nw=1.5E-07
XXI5 net0143 VDD VSS Q / INV pl=6E-08 pw=3.8E-07 nl=6E-08 nw=3E-07
XXI13 net0106 VDD VSS net24 / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI10 net0122 VDD VSS net0143 / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI4 CK VDD VSS net0106 / INV pl=6E-08 pw=2.1E-07 nl=6E-08 nw=1.7E-07
XXI9 net24 net0106 net46 net0122 VDD VSS / TG pl=6E-08 pw=1.9E-07 nl=6E-08
+ nw=1.5E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFSRX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFSRX0P5H7L CK D Q QN RN SN VDD VSS
*.PININFO CK:I D:I RN:I SN:I Q:O QN:O VDD:B VSS:B
MMN5 net062 SN VSS VSS nm1p2_lvt_lp W=240n L=60n m=1
MMN1 net093 CKN net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0144 net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN6 net093 R net062 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN4 net46 net33 net062 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMP4 net093 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP5 net54 R VDD VDD pm1p2_lvt_lp W=280n L=60n m=1
MMP2 net67 net0144 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net093 CKP net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=280n L=60n m=1
XXI29 net46 CKP CKN VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI30 D CKN CKP VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI3 net0144 VDD VSS Q / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI1 RN VDD VSS R / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI4 net093 VDD VSS QN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI0 CKN VDD VSS CKP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI2 net093 VDD VSS net0144 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI4 CK VDD VSS CKN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI9 CKP CKN net46 net093 VDD VSS / TG pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFSRX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFSRX1H7L CK D Q QN RN SN VDD VSS
*.PININFO CK:I D:I RN:I SN:I Q:O QN:O VDD:B VSS:B
MMN5 net062 SN VSS VSS nm1p2_lvt_lp W=240n L=60n m=1
MMN1 net093 CKN net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0144 net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN6 net093 R net062 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN4 net46 net33 net062 VSS nm1p2_lvt_lp W=215n L=60n m=1
MMP4 net093 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP5 net54 R VDD VDD pm1p2_lvt_lp W=300n L=60n m=1
MMP2 net67 net0144 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net093 CKP net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=300n L=60n m=1
XXI29 net46 CKP CKN VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI30 D CKN CKP VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI3 net0144 VDD VSS Q / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI1 RN VDD VSS R / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI5 net093 VDD VSS QN / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI0 CKN VDD VSS CKP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI2 net093 VDD VSS net0144 / INV pl=6E-08 pw=3E-07 nl=6E-08 nw=2.2E-07
XXI4 CK VDD VSS CKN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI9 CKP CKN net46 net093 VDD VSS / TG pl=6E-08 pw=3E-07 nl=6E-08 nw=2.2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFSRX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFSRX2H7L CK D Q QN RN SN VDD VSS
*.PININFO CK:I D:I RN:I SN:I Q:O QN:O VDD:B VSS:B
MMN5 net062 SN VSS VSS nm1p2_lvt_lp W=260n L=60n m=1
MMN1 net093 CKN net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0144 net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN6 net093 R net062 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN4 net46 net33 net062 VSS nm1p2_lvt_lp W=240n L=60n m=1
MMP4 net093 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP5 net54 R VDD VDD pm1p2_lvt_lp W=340n L=60n m=1
MMP2 net67 net0144 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net093 CKP net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=340n L=60n m=1
XXI29 net46 CKP CKN VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI30 D CKN CKP VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI3 net0144 VDD VSS Q / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI6 RN VDD VSS R / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI7 net093 VDD VSS QN / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI5 CKN VDD VSS CKP / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI8 net093 VDD VSS net0144 / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI4 CK VDD VSS CKN / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI9 CKP CKN net46 net093 VDD VSS / TG pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFSX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFSX0P5H7L CK D Q QN SN VDD VSS
*.PININFO CK:I D:I SN:I Q:O QN:O VDD:B VSS:B
MMN6 net056 SN VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMN1 net081 CKN net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0123 net056 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 net056 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMP0 net081 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP2 net67 net0123 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net081 CKP net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 VDD VDD pm1p2_lvt_lp W=280n L=60n m=1
XXI29 net46 CKP CKN VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI30 D CKN CKP VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI2 net0123 VDD VSS Q / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI3 net081 VDD VSS QN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI0 CKN VDD VSS CKP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI1 net081 VDD VSS net0123 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI4 CK VDD VSS CKN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI9 CKP CKN net46 net081 VDD VSS / TG pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFSX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFSX1H7L CK D Q QN SN VDD VSS
*.PININFO CK:I D:I SN:I Q:O QN:O VDD:B VSS:B
MMN6 net056 SN VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMN1 net081 CKN net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0123 net056 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 net056 VSS nm1p2_lvt_lp W=220n L=60n m=1
MMP0 net081 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP2 net67 net0123 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net081 CKP net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 VDD VDD pm1p2_lvt_lp W=300n L=60n m=1
XXI29 net46 CKP CKN VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI30 D CKN CKP VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI2 net0123 VDD VSS Q / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI5 net081 VDD VSS QN / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI0 CKN VDD VSS CKP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI1 net081 VDD VSS net0123 / INV pl=6E-08 pw=3E-07 nl=6E-08 nw=2.2E-07
XXI4 CK VDD VSS CKN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI9 CKP CKN net46 net081 VDD VSS / TG pl=6E-08 pw=3E-07 nl=6E-08 nw=2.2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFSX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFSX2H7L CK D Q QN SN VDD VSS
*.PININFO CK:I D:I SN:I Q:O QN:O VDD:B VSS:B
MMN6 net056 SN VSS VSS nm1p2_lvt_lp W=240n L=60n m=1
MMN1 net081 CKN net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0123 net056 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 net056 VSS nm1p2_lvt_lp W=240n L=60n m=1
MMP0 net081 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP2 net67 net0123 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net081 CKP net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 VDD VDD pm1p2_lvt_lp W=340n L=60n m=1
XXI29 net46 CKP CKN VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI30 D CKN CKP VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI6 net0123 VDD VSS Q / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI3 net081 VDD VSS QN / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI4 CKN VDD VSS CKP / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI5 net081 VDD VSS net0123 / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI4 CK VDD VSS CKN / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI9 CKP CKN net46 net081 VDD VSS / TG pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net15 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 net15 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP2 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFTRQX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFTRQX0P5H7L CK D Q RN VDD VSS
*.PININFO CK:I D:I RN:I Q:O VDD:B VSS:B
XXI17 D RN VDD VSS net030 / NAND2 pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2.4E-07
XXI18 net32 net24 net030 net33 VDD VSS / TG pl=6E-08 pw=2.8E-07 nl=6E-08
+ nw=2.4E-07
XXI14 net46 net24 net32 VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI9 net46 net24 net32 VDD VSS net25 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08
+ nw=2E-07
XXI15 net9 net32 net24 VDD VSS net25 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI7 net33 VDD VSS net46 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI13 net32 VDD VSS net24 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI12 net25 VDD VSS Q / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI10 net25 VDD VSS net9 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI4 CK VDD VSS net32 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net15 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 net15 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP2 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFTRQX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFTRQX1H7L CK D Q RN VDD VSS
*.PININFO CK:I D:I RN:I Q:O VDD:B VSS:B
XXI18 net32 net24 net034 net33 VDD VSS / TG pl=6E-08 pw=2.8E-07 nl=6E-08
+ nw=2.4E-07
XXI17 D RN VDD VSS net034 / NAND2 pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI14 net46 net24 net32 VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI9 net46 net24 net32 VDD VSS net25 / TSINV pl=6E-08 pw=3E-07 nl=6E-08
+ nw=2.2E-07
XXI15 net9 net32 net24 VDD VSS net25 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI7 net33 VDD VSS net46 / INV pl=6E-08 pw=3E-07 nl=6E-08 nw=2.2E-07
XXI13 net32 VDD VSS net24 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI12 net25 VDD VSS Q / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI10 net25 VDD VSS net9 / INV pl=6E-08 pw=3E-07 nl=6E-08 nw=2.2E-07
XXI4 CK VDD VSS net32 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net15 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 net15 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP2 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFTRQX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFTRQX2H7L CK D Q RN VDD VSS
*.PININFO CK:I D:I RN:I Q:O VDD:B VSS:B
XXI18 net32 net24 net034 net33 VDD VSS / TG pl=6E-08 pw=2.8E-07 nl=6E-08
+ nw=2.4E-07
XXI17 D RN VDD VSS net034 / NAND2 pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2.4E-07
XXI14 net46 net24 net32 VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI9 net46 net24 net32 VDD VSS net25 / TSINV pl=6E-08 pw=3.4E-07 nl=6E-08
+ nw=2.4E-07
XXI15 net9 net32 net24 VDD VSS net25 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XXI7 net33 VDD VSS net46 / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI13 net32 VDD VSS net24 / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI12 net25 VDD VSS Q / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XXI10 net25 VDD VSS net9 / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI4 CK VDD VSS net32 / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFX0P5H7L CK D Q QN VDD VSS
*.PININFO CK:I D:I Q:O QN:O VDD:B VSS:B
XI9 net9 CKN CKP VDD VSS net25 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08 nw=1.5E-07
XI10 net46 CKP CKN VDD VSS net25 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI11 net46 CKP CKN VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XI14 D CKN CKP VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI7 net9 VDD VSS QN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI16 net25 VDD VSS Q / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI8 CK VDD VSS CKN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI12 net33 VDD VSS net46 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI13 CKN VDD VSS CKP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI10 net25 VDD VSS net9 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFX1H7L CK D Q QN VDD VSS
*.PININFO CK:I D:I Q:O QN:O VDD:B VSS:B
XI2 net46 CKP CKN VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08 nw=1.5E-07
XXI6 D CKN CKP VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI3 net46 CKP CKN VDD VSS net25 / TSINV pl=6E-08 pw=3E-07 nl=6E-08 nw=2.2E-07
XI4 net9 CKN CKP VDD VSS net25 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08 nw=1.5E-07
XI1 net33 VDD VSS net46 / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI0 CKN VDD VSS CKP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI12 net25 VDD VSS Q / INV pl=6E-08 pw=3E-07 nl=6E-08 nw=2.4E-07
XXI10 net25 VDD VSS net9 / INV pl=6E-08 pw=3E-07 nl=6E-08 nw=2.2E-07
XI5 net9 VDD VSS QN / INV pl=6E-08 pw=3E-07 nl=6E-08 nw=2.4E-07
XXI4 CK VDD VSS CKN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFX2H7L CK D Q QN VDD VSS
*.PININFO CK:I D:I Q:O QN:O VDD:B VSS:B
XI7 net33 VDD VSS net46 / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI6 CKN VDD VSS CKP / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XXI12 net25 VDD VSS Q / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI8 net25 VDD VSS net9 / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI9 net9 VDD VSS QN / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XXI4 CK VDD VSS CKN / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI2 net46 CKP CKN VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08 nw=1.5E-07
XXI6 D CKN CKP VDD VSS net33 / TSINV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI3 net46 CKP CKN VDD VSS net25 / TSINV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI4 net9 CKN CKP VDD VSS net25 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08 nw=1.5E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DFFX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT DFFX3H7L CK D Q QN VDD VSS
*.PININFO CK:I D:I Q:O QN:O VDD:B VSS:B
XI13 net46 CKP CKN VDD VSS net33 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08
+ nw=1.5E-07
XI12 D CKN CKP VDD VSS net33 / TSINV pl=60n pw=340n nl=60n nw=240n
XI11 net46 CKP CKN VDD VSS net25 / TSINV pl=60n pw=360n nl=60n nw=260n
XI10 net9 CKN CKP VDD VSS net25 / TSINV pl=6E-08 pw=1.5E-07 nl=6E-08 nw=1.5E-07
XI19 net33 VDD VSS net46 / INV pl=60n pw=360n nl=60n nw=260n
XI18 CKN VDD VSS CKP / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI17 net25 VDD VSS Q / INV pl=60n pw=600n nl=60n nw=420n
XI16 net25 VDD VSS net9 / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI15 net9 VDD VSS QN / INV pl=60n pw=600n nl=60n nw=420n
XI14 CK VDD VSS CKN / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DLY1X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT DLY1X2H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XI3 net1 VDD VSS Y / INV pl=60n pw=380n nl=60n nw=190n
XI2 net2 VDD VSS net1 / INV pl=60n pw=270n nl=60n nw=150n
XI1 net3 VDD VSS net2 / INV pl=60n pw=190n nl=60n nw=150n
XI0 A VDD VSS net3 / INV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DLY1X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT DLY1X6H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XI0 A VDD VSS net013 / INV pl=60n pw=190n nl=60n nw=150n
XI1 net013 VDD VSS net014 / INV pl=60n pw=190n nl=60n nw=150n
XI2 net014 VDD VSS net015 / INV pl=60n pw=290n nl=60n nw=150n
XI3 net015 VDD VSS Y / INV pl=60n pw=1.14u nl=60n nw=570n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DLY2X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT DLY2X2H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XI3 net013 VDD VSS Y / INV pl=60n pw=380n nl=60n nw=190n
XI2 net014 VDD VSS net013 / INV pl=120n pw=230n nl=120n nw=150n
XI1 net015 VDD VSS net014 / INV pl=120n pw=190n nl=120n nw=150n
XI0 A VDD VSS net015 / INV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DLY2X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT DLY2X6H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XI0 A VDD VSS net013 / INV pl=60n pw=190n nl=60n nw=150n
XI1 net013 VDD VSS net014 / INV pl=120n pw=190n nl=120n nw=150n
XI2 net014 VDD VSS net015 / INV pl=120n pw=260n nl=120n nw=150n
XI3 net015 VDD VSS Y / INV pl=60n pw=1.14u nl=60n nw=570n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DLY3X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT DLY3X2H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XI0 A VDD VSS net013 / INV pl=60n pw=190n nl=60n nw=150n
XI1 net013 VDD VSS net014 / INV pl=180n pw=190n nl=180n nw=150n
XI2 net014 VDD VSS net015 / INV pl=180n pw=200n nl=180n nw=150n
XI3 net015 VDD VSS Y / INV pl=60n pw=380n nl=60n nw=190n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DLY3X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT DLY3X6H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XI3 net013 VDD VSS Y / INV pl=60n pw=1.14u nl=60n nw=570n
XI2 net014 VDD VSS net013 / INV pl=180n pw=250n nl=180n nw=160n
XI1 net015 VDD VSS net014 / INV pl=180n pw=190n nl=180n nw=150n
XI0 A VDD VSS net015 / INV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DLY4X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT DLY4X2H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XI3 net013 VDD VSS Y / INV pl=60n pw=380n nl=60n nw=190n
XI2 net014 VDD VSS net013 / INV pl=240n pw=190n nl=240n nw=150n
XI1 net015 VDD VSS net014 / INV pl=240n pw=190n nl=240n nw=150n
XI0 A VDD VSS net015 / INV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    DLY4X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT DLY4X6H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XI0 A VDD VSS net013 / INV pl=60n pw=190n nl=60n nw=150n
XI1 net013 VDD VSS net014 / INV pl=240n pw=190n nl=240n nw=150n
XI2 net014 VDD VSS net015 / INV pl=240n pw=220n nl=240n nw=150n
XI3 net015 VDD VSS Y / INV pl=60n pw=1.14u nl=60n nw=570n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    EDFFQX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT EDFFQX0P5H7L CK D E Q VDD VSS
*.PININFO CK:I D:I E:I Q:O VDD:B VSS:B
XXI18 net32 net24 net030 net33 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
XXI14 net46 net24 net32 VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI17 D E net057 VDD VSS net030 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI19 net9 net057 E VDD VSS net030 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI9 net46 net24 net32 VDD VSS net25 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI15 net9 net32 net24 VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI20 E VDD VSS net057 / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=280n nl=60n nw=200n
XXI13 net32 VDD VSS net24 / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net25 VDD VSS Q / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XXI4 CK VDD VSS net32 / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    EDFFQX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT EDFFQX1H7L CK D E Q VDD VSS
*.PININFO CK:I D:I E:I Q:O VDD:B VSS:B
XXI18 net32 net24 net030 net33 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
XXI14 net46 net24 net32 VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI17 D E net057 VDD VSS net030 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI19 net9 net057 E VDD VSS net030 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI9 net46 net24 net32 VDD VSS net25 / TSINV pl=60n pw=300n nl=60n nw=220n
XXI15 net9 net32 net24 VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI20 E VDD VSS net057 / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=280n nl=60n nw=200n
XXI13 net32 VDD VSS net24 / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net25 VDD VSS Q / INV pl=60n pw=340n nl=60n nw=240n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XXI4 CK VDD VSS net32 / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    EDFFQX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT EDFFQX2H7L CK D E Q VDD VSS
*.PININFO CK:I D:I E:I Q:O VDD:B VSS:B
XXI18 net32 net24 net030 net33 VDD VSS / TG pl=60n pw=340n nl=60n nw=240n
XXI14 net46 net24 net32 VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI17 D E net057 VDD VSS net030 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI19 net9 net057 E VDD VSS net030 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI9 net46 net24 net32 VDD VSS net25 / TSINV pl=60n pw=340n nl=60n nw=240n
XXI15 net9 net32 net24 VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI20 E VDD VSS net057 / INV pl=60n pw=340n nl=60n nw=240n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=280n nl=60n nw=200n
XXI13 net32 VDD VSS net24 / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net25 VDD VSS Q / INV pl=60n pw=400n nl=60n nw=280n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XXI4 CK VDD VSS net32 / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    ESDFFQX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT ESDFFQX0P5H7L CK D E Q SE SI VDD VSS
*.PININFO CK:I D:I E:I SE:I SI:I Q:O VDD:B VSS:B
XXI21 c cn net46 net25 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
XXI20 SEN SE net034 net046 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
XI2 net046 cn c VDD VSS net33 / TSINV pl=60n pw=300n nl=60n nw=220n
XXI25 net9 EN E VDD VSS net034 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI24 D E EN VDD VSS net034 / TSINV pl=60n pw=300n nl=60n nw=220n
XXI14 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI22 SI SE SEN VDD VSS net046 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI15 net9 cn c VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI26 E VDD VSS EN / INV pl=60n pw=280n nl=60n nw=200n
XXI23 SE VDD VSS SEN / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=280n nl=60n nw=200n
XXI13 cn VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net25 VDD VSS Q / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XXI4 CK VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    ESDFFQX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT ESDFFQX1H7L CK D E Q SE SI VDD VSS
*.PININFO CK:I D:I E:I SE:I SI:I Q:O VDD:B VSS:B
XXI21 c cn net46 net25 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
XXI20 SEN SE net034 net046 VDD VSS / TG pl=60n pw=320n nl=60n nw=240n
XXI25 net9 EN E VDD VSS net034 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI24 D E EN VDD VSS net034 / TSINV pl=60n pw=320n nl=60n nw=240n
XXI14 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI22 SI SE SEN VDD VSS net046 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI19 net046 cn c VDD VSS net33 / TSINV pl=60n pw=320n nl=60n nw=240n
XXI15 net9 cn c VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI26 E VDD VSS EN / INV pl=60n pw=280n nl=60n nw=200n
XXI23 SE VDD VSS SEN / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=300n nl=60n nw=220n
XXI13 cn VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net25 VDD VSS Q / INV pl=60n pw=340n nl=60n nw=240n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XXI4 CK VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    ESDFFQX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT ESDFFQX2H7L CK D E Q SE SI VDD VSS
*.PININFO CK:I D:I E:I SE:I SI:I Q:O VDD:B VSS:B
XXI20 SEN SE net034 net046 VDD VSS / TG pl=60n pw=320n nl=60n nw=240n
XXI21 c cn net46 net25 VDD VSS / TG pl=60n pw=340n nl=60n nw=240n
XXI15 net9 cn c VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI19 net046 cn c VDD VSS net33 / TSINV pl=60n pw=320n nl=60n nw=240n
XXI22 SI SE SEN VDD VSS net046 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI14 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI24 D E EN VDD VSS net034 / TSINV pl=60n pw=320n nl=60n nw=240n
XXI25 net9 EN E VDD VSS net034 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI4 CK VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net25 VDD VSS Q / INV pl=60n pw=400n nl=60n nw=280n
XXI13 cn VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=340n nl=60n nw=240n
XXI23 SE VDD VSS SEN / INV pl=60n pw=280n nl=60n nw=200n
XXI26 E VDD VSS EN / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    FILLCAP16H7L
* View Name:    schematic
************************************************************************

.SUBCKT FILLCAP16H7L VDD VSS
*.PININFO VDD:B VSS:B
MMM1 net5 net7 VSS VSS nm1p2_lvt_lp W=200n L=2.78u m=1
MMM0 net7 net5 VDD VDD pm1p2_lvt_lp W=300n L=2.78u m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    FILLCAP32H7L
* View Name:    schematic
************************************************************************

.SUBCKT FILLCAP32H7L VDD VSS
*.PININFO VDD:B VSS:B
MMM1 net5 net7 VSS VSS nm1p2_lvt_lp W=200n L=5.98u m=1
MMM0 net7 net5 VDD VDD pm1p2_lvt_lp W=300n L=5.98u m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    FILLCAP4H7L
* View Name:    schematic
************************************************************************

.SUBCKT FILLCAP4H7L VDD VSS
*.PININFO VDD:B VSS:B
MMM1 net1 net3 VSS VSS nm1p2_lvt_lp W=200n L=380n m=1
MMM0 net3 net1 VDD VDD pm1p2_lvt_lp W=300n L=380n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    FILLCAP8H7L
* View Name:    schematic
************************************************************************

.SUBCKT FILLCAP8H7L VDD VSS
*.PININFO VDD:B VSS:B
MMM0 net7 net5 VDD VDD pm1p2_lvt_lp W=300n L=1.18u m=1
MMM1 net5 net7 VSS VSS nm1p2_lvt_lp W=200n L=1.18u m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    FILLER16H7L
* View Name:    schematic
************************************************************************

.SUBCKT FILLER16H7L VDD VSS
*.PININFO VDD:B VSS:B
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    FILLER1H7L
* View Name:    schematic
************************************************************************

.SUBCKT FILLER1H7L VDD VSS
*.PININFO VDD:B VSS:B
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    FILLER2H7L
* View Name:    schematic
************************************************************************

.SUBCKT FILLER2H7L VDD VSS
*.PININFO VDD:B VSS:B
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    FILLER32H7L
* View Name:    schematic
************************************************************************

.SUBCKT FILLER32H7L VDD VSS
*.PININFO VDD:B VSS:B
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    FILLER4H7L
* View Name:    schematic
************************************************************************

.SUBCKT FILLER4H7L VDD VSS
*.PININFO VDD:B VSS:B
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    FILLER64H7L
* View Name:    schematic
************************************************************************

.SUBCKT FILLER64H7L VDD VSS
*.PININFO VDD:B VSS:B
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    FILLER8H7L
* View Name:    schematic
************************************************************************

.SUBCKT FILLER8H7L VDD VSS
*.PININFO VDD:B VSS:B
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    FILLTAPH7L
* View Name:    schematic
************************************************************************

.SUBCKT FILLTAPH7L VDD VSS
*.PININFO VDD:I VSS:I
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NOR2
* View Name:    schematic
************************************************************************

.SUBCKT NOR2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 Y A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 Y B net018 VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP2 net018 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    ICGNX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT ICGNX0P5H7L CKN E ECK VDD VSS
*.PININFO CKN:I E:I ECK:O VDD:B VSS:B
XXI1 net9 CKN VDD VSS net14 / NOR2 pl=60n pw=320n nl=60n nw=200n
XXI6 CKN VDD VSS net8 / INV pl=60n pw=280n nl=60n nw=200n
XXI5 net8 VDD VSS net11 / INV pl=60n pw=280n nl=60n nw=200n
XXI2 net9 VDD VSS net6 / INV pl=60n pw=280n nl=60n nw=200n
XXI0 net14 VDD VSS ECK / INV pl=60n pw=280n nl=60n nw=200n
XXI4 net6 net8 net11 VDD VSS net9 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI3 E net11 net8 VDD VSS net9 / TSINV pl=60n pw=320n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NOR2
* View Name:    schematic
************************************************************************

.SUBCKT NOR2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 Y A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 Y B net018 VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP2 net018 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    ICGNX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT ICGNX1H7L CKN E ECK VDD VSS
*.PININFO CKN:I E:I ECK:O VDD:B VSS:B
XXI1 net9 CKN VDD VSS net14 / NOR2 pl=60n pw=320n nl=60n nw=200n
XXI6 CKN VDD VSS net8 / INV pl=60n pw=280n nl=60n nw=200n
XXI5 net8 VDD VSS net11 / INV pl=60n pw=280n nl=60n nw=200n
XXI2 net9 VDD VSS net6 / INV pl=60n pw=280n nl=60n nw=200n
XXI0 net14 VDD VSS ECK / INV pl=60n pw=340n nl=60n nw=240n
XXI4 net6 net8 net11 VDD VSS net9 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI3 E net11 net8 VDD VSS net9 / TSINV pl=60n pw=320n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NOR2
* View Name:    schematic
************************************************************************

.SUBCKT NOR2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 Y A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 Y B net018 VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP2 net018 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    ICGNX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT ICGNX2H7L CKN E ECK VDD VSS
*.PININFO CKN:I E:I ECK:O VDD:B VSS:B
XXI1 net9 CKN VDD VSS net14 / NOR2 pl=60n pw=320n nl=60n nw=200n
XXI6 CKN VDD VSS net8 / INV pl=60n pw=280n nl=60n nw=200n
XXI5 net8 VDD VSS net11 / INV pl=60n pw=280n nl=60n nw=200n
XXI2 net9 VDD VSS net6 / INV pl=60n pw=280n nl=60n nw=200n
XXI0 net14 VDD VSS ECK / INV pl=60n pw=400n nl=60n nw=280n
XXI4 net6 net8 net11 VDD VSS net9 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI3 E net11 net8 VDD VSS net9 / TSINV pl=60n pw=320n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NOR2
* View Name:    schematic
************************************************************************

.SUBCKT NOR2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 Y A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 Y B net018 VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP2 net018 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    ICGNX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT ICGNX3H7L CKN E ECK VDD VSS
*.PININFO CKN:I E:I ECK:O VDD:B VSS:B
XXI1 net9 CKN VDD VSS net14 / NOR2 pl=60n pw=360n nl=60n nw=220n
XXI6 CKN VDD VSS net8 / INV pl=60n pw=280n nl=60n nw=200n
XXI5 net8 VDD VSS net11 / INV pl=60n pw=280n nl=60n nw=200n
XXI2 net9 VDD VSS net6 / INV pl=60n pw=280n nl=60n nw=200n
XXI0 net14 VDD VSS ECK / INV pl=60n pw=600n nl=60n nw=420n
XXI4 net6 net8 net11 VDD VSS net9 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI3 E net11 net8 VDD VSS net9 / TSINV pl=60n pw=320n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NOR2
* View Name:    schematic
************************************************************************

.SUBCKT NOR2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 Y A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 Y B net018 VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP2 net018 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    ICGNX4H7L
* View Name:    schematic
************************************************************************

.SUBCKT ICGNX4H7L CKN E ECK VDD VSS
*.PININFO CKN:I E:I ECK:O VDD:B VSS:B
XXI1 net9 CKN VDD VSS net14 / NOR2 pl=60n pw=360n nl=60n nw=220n
XXI6 CKN VDD VSS net8 / INV pl=60n pw=280n nl=60n nw=200n
XXI5 net8 VDD VSS net11 / INV pl=60n pw=280n nl=60n nw=200n
XXI2 net9 VDD VSS net6 / INV pl=60n pw=280n nl=60n nw=200n
XXI0 net14 VDD VSS ECK / INV pl=60n pw=800n nl=60n nw=560n
XXI4 net6 net8 net11 VDD VSS net9 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI3 E net11 net8 VDD VSS net9 / TSINV pl=60n pw=320n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net15 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 net15 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP2 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    ICGX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT ICGX0P5H7L CK E ECK VDD VSS
*.PININFO CK:I E:I ECK:O VDD:B VSS:B
XXI1 net6 CK VDD VSS net14 / NAND2 pl=60n pw=200n nl=60n nw=200n
XXI6 CK VDD VSS net8 / INV pl=60n pw=280n nl=60n nw=200n
XXI5 net8 VDD VSS net11 / INV pl=60n pw=280n nl=60n nw=200n
XXI2 net9 VDD VSS net6 / INV pl=60n pw=280n nl=60n nw=200n
XXI0 net14 VDD VSS ECK / INV pl=60n pw=280n nl=60n nw=200n
XXI4 net6 net11 net8 VDD VSS net9 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI3 E net8 net11 VDD VSS net9 / TSINV pl=60n pw=320n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net15 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 net15 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP2 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    ICGX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT ICGX1H7L CK E ECK VDD VSS
*.PININFO CK:I E:I ECK:O VDD:B VSS:B
XXI1 net6 CK VDD VSS net14 / NAND2 pl=60n pw=200n nl=60n nw=220n
XXI6 CK VDD VSS net8 / INV pl=60n pw=280n nl=60n nw=200n
XXI5 net8 VDD VSS net11 / INV pl=60n pw=280n nl=60n nw=200n
XXI2 net9 VDD VSS net6 / INV pl=60n pw=280n nl=60n nw=200n
XXI0 net14 VDD VSS ECK / INV pl=60n pw=340n nl=60n nw=240n
XXI4 net6 net11 net8 VDD VSS net9 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI3 E net8 net11 VDD VSS net9 / TSINV pl=60n pw=320n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net15 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 net15 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP2 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    ICGX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT ICGX2H7L CK E ECK VDD VSS
*.PININFO CK:I E:I ECK:O VDD:B VSS:B
XXI1 net6 CK VDD VSS net14 / NAND2 pl=60n pw=200n nl=60n nw=220n
XXI6 CK VDD VSS net8 / INV pl=60n pw=280n nl=60n nw=200n
XXI2 net9 VDD VSS net6 / INV pl=60n pw=280n nl=60n nw=200n
XXI5 net8 VDD VSS net11 / INV pl=60n pw=280n nl=60n nw=200n
XXI0 net14 VDD VSS ECK / INV pl=60n pw=400n nl=60n nw=280n
XXI3 E net8 net11 VDD VSS net9 / TSINV pl=60n pw=320n nl=60n nw=200n
XXI4 net6 net11 net8 VDD VSS net9 / TSINV pl=60n pw=150n nl=60n nw=150n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net15 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 net15 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP2 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    ICGX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT ICGX3H7L CK E ECK VDD VSS
*.PININFO CK:I E:I ECK:O VDD:B VSS:B
XXI1 net6 CK VDD VSS net14 / NAND2 pl=60n pw=200n nl=60n nw=280n
XXI6 CK VDD VSS net8 / INV pl=60n pw=280n nl=60n nw=200n
XXI2 net9 VDD VSS net6 / INV pl=60n pw=280n nl=60n nw=200n
XXI5 net8 VDD VSS net11 / INV pl=60n pw=280n nl=60n nw=200n
XXI0 net14 VDD VSS ECK / INV pl=60n pw=600n nl=60n nw=420n
XXI3 E net8 net11 VDD VSS net9 / TSINV pl=60n pw=320n nl=60n nw=200n
XXI4 net6 net11 net8 VDD VSS net9 / TSINV pl=60n pw=150n nl=60n nw=150n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net15 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 net15 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP2 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    ICGX4H7L
* View Name:    schematic
************************************************************************

.SUBCKT ICGX4H7L CK E ECK VDD VSS
*.PININFO CK:I E:I ECK:O VDD:B VSS:B
XXI1 net6 CK VDD VSS net14 / NAND2 pl=60n pw=200n nl=60n nw=280n
XXI6 CK VDD VSS net8 / INV pl=60n pw=280n nl=60n nw=200n
XXI5 net8 VDD VSS net11 / INV pl=60n pw=280n nl=60n nw=200n
XXI2 net9 VDD VSS net6 / INV pl=60n pw=280n nl=60n nw=200n
XXI0 net14 VDD VSS ECK / INV pl=60n pw=800n nl=60n nw=560n
XXI4 net6 net11 net8 VDD VSS net9 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI3 E net8 net11 VDD VSS net9 / TSINV pl=60n pw=320n nl=60n nw=200n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    INVX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT INVX0P5H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI0 A VDD VSS Y / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    INVX0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT INVX0P7H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI0 A VDD VSS Y / INV pl=6e-08 pw=2.22e-07 nl=6e-08 nw=1.74e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    INVX10H7L
* View Name:    schematic
************************************************************************

.SUBCKT INVX10H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI0 A VDD VSS Y / INV pl=6e-08 pw=1.9e-06 nl=6e-08 nw=1.5e-06
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    INVX12H7L
* View Name:    schematic
************************************************************************

.SUBCKT INVX12H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI0 A VDD VSS Y / INV pl=6e-08 pw=2.28e-06 nl=6e-08 nw=1.8e-06
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    INVX16H7L
* View Name:    schematic
************************************************************************

.SUBCKT INVX16H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI0 A VDD VSS Y / INV pl=6e-08 pw=3.04e-06 nl=6e-08 nw=2.4e-06
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    INVX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT INVX1H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI0 A VDD VSS Y / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    INVX1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT INVX1P4H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI0 A VDD VSS Y / INV pl=6e-08 pw=3.14e-07 nl=6e-08 nw=2.46e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    INVX20H7L
* View Name:    schematic
************************************************************************

.SUBCKT INVX20H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI0 A VDD VSS Y / INV pl=6e-08 pw=3.8e-06 nl=6e-08 nw=3e-06
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    INVX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT INVX2H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI0 A VDD VSS Y / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    INVX2P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT INVX2P5H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI0 A VDD VSS Y / INV pl=6e-08 pw=4.75e-07 nl=6e-08 nw=3.75e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    INVX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT INVX3H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI0 A VDD VSS Y / INV pl=6e-08 pw=5.7e-07 nl=6e-08 nw=4.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    INVX3P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT INVX3P5H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI0 A VDD VSS Y / INV pl=6e-08 pw=6.65e-07 nl=6e-08 nw=5.25e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    INVX4H7L
* View Name:    schematic
************************************************************************

.SUBCKT INVX4H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI0 A VDD VSS Y / INV pl=6e-08 pw=7.6e-07 nl=6e-08 nw=6e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    INVX5H7L
* View Name:    schematic
************************************************************************

.SUBCKT INVX5H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI0 A VDD VSS Y / INV pl=6e-08 pw=9.5e-07 nl=6e-08 nw=7.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    INVX6H7L
* View Name:    schematic
************************************************************************

.SUBCKT INVX6H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI0 A VDD VSS Y / INV pl=6e-08 pw=1.14e-06 nl=6e-08 nw=9e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    INVX7H7L
* View Name:    schematic
************************************************************************

.SUBCKT INVX7H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI0 A VDD VSS Y / INV pl=6e-08 pw=1.33e-06 nl=6e-08 nw=1.05e-06
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    INVX8H7L
* View Name:    schematic
************************************************************************

.SUBCKT INVX8H7L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
XXI0 A VDD VSS Y / INV pl=6e-08 pw=1.52e-06 nl=6e-08 nw=1.2e-06
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATHRX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATHRX0P5H7L D G Q QN RN VDD VSS
*.PININFO D:I G:I RN:I Q:O QN:O VDD:B VSS:B
MMN3 net44 RN VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN2 net47 D net44 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN4 net41 netqn net38 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net38 RN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 netq GN net41 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP1 net47 D VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP4 netq GP net059 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP5 net059 netqn VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 netq RN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
XI4 netq VDD VSS Q / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI2 netq VDD VSS netqn / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI3 netqn VDD VSS QN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI1 GN VDD VSS GP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI0 G VDD VSS GN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI9 GP GN net47 netq VDD VSS / TG pl=6E-08 pw=2.7E-07 nl=6E-08 nw=1.95E-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATHRX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATHRX1H7L D G Q QN RN VDD VSS
*.PININFO D:I G:I RN:I Q:O QN:O VDD:B VSS:B
MNM0 net44 RN VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN2 net47 D net44 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN4 net41 netqn net38 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net38 RN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 netq GN net41 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP1 net47 D VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP4 netq GP net059 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP5 net059 netqn VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 netq RN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
XI4 netq VDD VSS Q / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI8 netq VDD VSS netqn / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI7 netqn VDD VSS QN / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI6 GN VDD VSS GP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI0 G VDD VSS GN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XXI9 GP GN net47 netq VDD VSS / TG pl=6E-08 pw=2.7E-07 nl=6E-08 nw=1.95E-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATHRX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATHRX2H7L D G Q QN RN VDD VSS
*.PININFO D:I G:I RN:I Q:O QN:O VDD:B VSS:B
MNM0 net47 D net44 VSS nm1p2_lvt_lp W=240n L=60n m=1
MMN3 net44 RN VSS VSS nm1p2_lvt_lp W=240n L=60n m=1
MMN4 net41 netqn net38 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net38 RN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 netq GN net41 VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM0 net47 D VDD VDD pm1p2_lvt_lp W=340n L=60n m=1
MMP4 netq GP net059 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP5 net059 netqn VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 netq RN VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
XI6 GN VDD VSS GP / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI10 netqn VDD VSS QN / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI9 netq VDD VSS netqn / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI4 netq VDD VSS Q / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI5 G VDD VSS GN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI7 GP GN net47 netq VDD VSS / TG pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATHSRX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATHSRX0P5H7L D G Q QN RN SN VDD VSS
*.PININFO D:I G:I RN:I SN:I Q:O QN:O VDD:B VSS:B
MNM1 net47 D net44 VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM2 net41 netqn net44 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM3 net0154 GN net41 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net0154 S VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM4 net44 RN VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MPM2 net052 netqn net058 VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM1 net0154 GP net052 VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM3 net47 D net058 VDD pm1p2_lvt_lp W=280n L=60n m=1
MPM0 net0154 RN net058 VDD pm1p2_lvt_lp W=200n L=60n m=1
MPM4 net058 S VDD VDD pm1p2_lvt_lp W=280n L=60n m=1
XI3 G VDD VSS GN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI0 GN VDD VSS GP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI2 net0154 VDD VSS netqn / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI5 net0154 VDD VSS Q / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI4 netqn VDD VSS QN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI1 SN VDD VSS S / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI7 GP GN net47 net0154 VDD VSS / TG pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATHSRX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATHSRX1H7L D G Q QN RN SN VDD VSS
*.PININFO D:I G:I RN:I SN:I Q:O QN:O VDD:B VSS:B
MNM1 net47 D net44 VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM2 net41 netqn net44 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM3 net0154 GN net41 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net0154 S VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM4 net44 RN VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MPM2 net052 netqn net058 VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM1 net0154 GP net052 VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM3 net47 D net058 VDD pm1p2_lvt_lp W=280n L=60n m=1
MPM0 net0154 RN net058 VDD pm1p2_lvt_lp W=200n L=60n m=1
MPM4 net058 S VDD VDD pm1p2_lvt_lp W=280n L=60n m=1
XI3 G VDD VSS GN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI0 GN VDD VSS GP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI2 net0154 VDD VSS netqn / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI6 net0154 VDD VSS Q / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI4 netqn VDD VSS QN / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI1 SN VDD VSS S / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI7 GP GN net47 net0154 VDD VSS / TG pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATHSRX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATHSRX2H7L D G Q QN RN SN VDD VSS
*.PININFO D:I G:I RN:I SN:I Q:O QN:O VDD:B VSS:B
MNM1 net47 D net44 VSS nm1p2_lvt_lp W=240n L=60n m=1
MNM2 net41 netqn net44 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM3 net0154 GN net41 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net0154 S VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM4 net44 RN VSS VSS nm1p2_lvt_lp W=240n L=60n m=1
MPM2 net052 netqn net058 VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM1 net0154 GP net052 VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM3 net47 D net058 VDD pm1p2_lvt_lp W=340n L=60n m=1
MPM0 net0154 RN net058 VDD pm1p2_lvt_lp W=200n L=60n m=1
MPM4 net058 S VDD VDD pm1p2_lvt_lp W=340n L=60n m=1
XI3 G VDD VSS GN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI2 net0154 VDD VSS netqn / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI8 net0154 VDD VSS Q / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI4 netqn VDD VSS QN / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI1 SN VDD VSS S / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI6 GN VDD VSS GP / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI7 GP GN net47 net0154 VDD VSS / TG pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATHSX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATHSX0P5H7L D G Q QN SN VDD VSS
*.PININFO D:I G:I SN:I Q:O QN:O VDD:B VSS:B
MNM1 net44 D VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM2 netq S VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN1 netq GN net38 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net38 netqn VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM2 net44 D net062 VDD pm1p2_lvt_lp W=320n L=60n m=1
MPM1 net065 S VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM0 net056 netqn net065 VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM3 net062 S VDD VDD pm1p2_lvt_lp W=320n L=60n m=1
MMP4 netq GP net056 VDD pm1p2_lvt_lp W=150n L=60n m=1
XI5 SN VDD VSS S / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI3 G VDD VSS GN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI0 netq VDD VSS Q / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI2 netq VDD VSS netqn / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI1 netqn VDD VSS QN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI4 GN VDD VSS GP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI7 GP GN net44 netq VDD VSS / TG pl=6E-08 pw=3.2E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATHSX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATHSX1H7L D G Q QN SN VDD VSS
*.PININFO D:I G:I SN:I Q:O QN:O VDD:B VSS:B
MNM1 net44 D VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM2 netq S VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN1 netq GN net38 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net38 netqn VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM2 net44 D net062 VDD pm1p2_lvt_lp W=320n L=60n m=1
MPM1 net065 S VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM0 net056 netqn net065 VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM4 net062 S VDD VDD pm1p2_lvt_lp W=320n L=60n m=1
MMP4 netq GP net056 VDD pm1p2_lvt_lp W=150n L=60n m=1
XI10 GN VDD VSS GP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI3 G VDD VSS GN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI0 netq VDD VSS Q / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI12 netq VDD VSS netqn / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI13 netqn VDD VSS QN / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI11 SN VDD VSS S / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI7 GP GN net44 netq VDD VSS / TG pl=6E-08 pw=3.2E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATHSX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATHSX2H7L D G Q QN SN VDD VSS
*.PININFO D:I G:I SN:I Q:O QN:O VDD:B VSS:B
MNM1 net44 D VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM2 netq S VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN1 netq GN net38 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net38 netqn VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM2 net44 D net062 VDD pm1p2_lvt_lp W=320n L=60n m=1
MPM1 net065 S VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM0 net056 netqn net065 VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM4 net062 S VDD VDD pm1p2_lvt_lp W=320n L=60n m=1
MMP4 netq GP net056 VDD pm1p2_lvt_lp W=150n L=60n m=1
XI11 SN VDD VSS S / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI15 netq VDD VSS Q / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI12 netq VDD VSS netqn / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI13 netqn VDD VSS QN / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI14 GN VDD VSS GP / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI3 G VDD VSS GN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI7 GP GN net44 netq VDD VSS / TG pl=6E-08 pw=3.2E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATHX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATHX0P5H7L D G Q QN VDD VSS
*.PININFO D:I G:I Q:O QN:O VDD:B VSS:B
XXI6 D GP GN VDD VSS net25 / TSINV pl=6e-08 pw=2.8e-07 nl=6e-08 nw=2e-07
XXI15 net9 GN GP VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI4 G VDD VSS GN / INV pl=60n pw=280n nl=60n nw=200n
XI2 net9 VDD VSS QN / INV pl=60n pw=280n nl=60n nw=200n
XXI13 GN VDD VSS GP / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XI3 net25 VDD VSS Q / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATHX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATHX1H7L D G Q QN VDD VSS
*.PININFO D:I G:I Q:O QN:O VDD:B VSS:B
XI9 D GP GN VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI15 net9 GN GP VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI4 G VDD VSS GN / INV pl=60n pw=280n nl=60n nw=200n
XI8 GN VDD VSS GP / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XI0 net25 VDD VSS Q / INV pl=60n pw=340n nl=60n nw=240n
XI1 net9 VDD VSS QN / INV pl=60n pw=340n nl=60n nw=240n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATHX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATHX2H7L D G Q QN VDD VSS
*.PININFO D:I G:I Q:O QN:O VDD:B VSS:B
XXI6 D GP GN VDD VSS net25 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI15 net9 GN GP VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XI11 GN VDD VSS GP / INV pl=60n pw=280n nl=60n nw=200n
XI9 G VDD VSS GN / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XI2 net25 VDD VSS Q / INV pl=60n pw=400n nl=60n nw=280n
XI1 net9 VDD VSS QN / INV pl=60n pw=400n nl=60n nw=280n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATHX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATHX3H7L D G Q QN VDD VSS
*.PININFO D:I G:I Q:O QN:O VDD:B VSS:B
XXI6 D GP GN VDD VSS net25 / TSINV pl=6e-08 pw=3.4e-07 nl=6e-08 nw=2.4e-07
XXI15 net9 GN GP VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI4 G VDD VSS GN / INV pl=60n pw=280n nl=60n nw=200n
XXI13 GN VDD VSS GP / INV pl=60n pw=340n nl=60n nw=240n
XXI7 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XI4 net25 VDD VSS Q / INV pl=60n pw=600n nl=60n nw=420n
XI1 net9 VDD VSS QN / INV pl=60n pw=600n nl=60n nw=420n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATHX4H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATHX4H7L D G Q QN VDD VSS
*.PININFO D:I G:I Q:O QN:O VDD:B VSS:B
XXI6 D GP GN VDD VSS net25 / TSINV pl=6e-08 pw=3.4e-07 nl=6e-08 nw=2.4e-07
XXI15 net9 GN GP VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI4 G VDD VSS GN / INV pl=60n pw=280n nl=60n nw=200n
XXI13 GN VDD VSS GP / INV pl=60n pw=340n nl=60n nw=240n
XXI7 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XI3 net25 VDD VSS Q / INV pl=60n pw=800n nl=60n nw=560n
XI1 net9 VDD VSS QN / INV pl=60n pw=800n nl=60n nw=560n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATLRX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATLRX0P5H7L D GN Q QN RN VDD VSS
*.PININFO D:I GN:I RN:I Q:O QN:O VDD:B VSS:B
MNM4 net47 D net12 VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM3 net12 RN VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM2 netq GB net52 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net52 netqn net51 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net51 RN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM3 netq RN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MPM2 net47 D VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM1 net53 netqn VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM0 netq GP net53 VDD pm1p2_lvt_lp W=150n L=60n m=1
XI1 GP VDD VSS GB / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI0 GN VDD VSS GP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI2 netq VDD VSS netqn / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI3 netqn VDD VSS QN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI5 netq VDD VSS Q / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI4 GP GB net47 netq VDD VSS / TG pl=6E-08 pw=2.7E-07 nl=6E-08 nw=1.95E-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATLRX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATLRX1H7L D GN Q QN RN VDD VSS
*.PININFO D:I GN:I RN:I Q:O QN:O VDD:B VSS:B
MNM4 net47 D net29 VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM3 net29 RN VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM2 netq GB net66 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net66 netqn net67 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net67 RN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM3 netq RN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MPM2 net47 D VDD VDD pm1p2_lvt_lp W=280n L=60n m=1
MPM1 net65 netqn VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM0 netq GP net65 VDD pm1p2_lvt_lp W=150n L=60n m=1
XI11 GP VDD VSS GB / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI12 GN VDD VSS GP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI13 netq VDD VSS netqn / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI14 netqn VDD VSS QN / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI16 netq VDD VSS Q / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI15 GP GB net47 netq VDD VSS / TG pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATLRX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATLRX2H7L D GN Q QN RN VDD VSS
*.PININFO D:I GN:I RN:I Q:O QN:O VDD:B VSS:B
MNM4 net47 D net29 VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM3 net29 RN VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM2 netq GB net66 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net66 netqn net67 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net67 RN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM3 netq RN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MPM2 net47 D VDD VDD pm1p2_lvt_lp W=280n L=60n m=1
MPM1 net65 netqn VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM0 netq GP net65 VDD pm1p2_lvt_lp W=150n L=60n m=1
XI11 GP VDD VSS GB / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI12 GN VDD VSS GP / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI13 netq VDD VSS netqn / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI14 netqn VDD VSS QN / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI16 netq VDD VSS Q / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI15 GP GB net47 netq VDD VSS / TG pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATLSRX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATLSRX0P5H7L D GN Q QN RN SN VDD VSS
*.PININFO D:I GN:I RN:I SN:I Q:O QN:O VDD:B VSS:B
XI3 GN VDD VSS G / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI0 G VDD VSS GB / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI2 net0102 VDD VSS netqn / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI4 netqn VDD VSS QN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI5 net0102 VDD VSS Q / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI1 SN VDD VSS S / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
MNM3 net0102 GB net41 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net0102 S VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM1 net47 D net44 VSS nm1p2_lvt_lp W=240n L=60n m=1
MNM2 net41 netqn net44 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM4 net44 RN VSS VSS nm1p2_lvt_lp W=240n L=60n m=1
XI7 G GB net47 net0102 VDD VSS / TG pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
MPM4 net059 S VDD VDD pm1p2_lvt_lp W=340n L=60n m=1
MPM2 net053 netqn net059 VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM3 net47 D net059 VDD pm1p2_lvt_lp W=340n L=60n m=1
MPM0 net0102 RN net059 VDD pm1p2_lvt_lp W=200n L=60n m=1
MPM1 net0102 G net053 VDD pm1p2_lvt_lp W=150n L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATLSRX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATLSRX1H7L D GN Q QN RN SN VDD VSS
*.PININFO D:I GN:I RN:I SN:I Q:O QN:O VDD:B VSS:B
XI3 GN VDD VSS G / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI0 G VDD VSS GB / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI2 net0102 VDD VSS netqn / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI4 netqn VDD VSS QN / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI5 net0102 VDD VSS Q / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI1 SN VDD VSS S / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
MNM3 net0102 GB net41 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net0102 S VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM1 net47 D net44 VSS nm1p2_lvt_lp W=240n L=60n m=1
MNM2 net41 netqn net44 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM4 net44 RN VSS VSS nm1p2_lvt_lp W=240n L=60n m=1
XI7 G GB net47 net0102 VDD VSS / TG pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
MPM4 net059 S VDD VDD pm1p2_lvt_lp W=340n L=60n m=1
MPM2 net053 netqn net059 VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM3 net47 D net059 VDD pm1p2_lvt_lp W=340n L=60n m=1
MPM0 net0102 RN net059 VDD pm1p2_lvt_lp W=200n L=60n m=1
MPM1 net0102 G net053 VDD pm1p2_lvt_lp W=150n L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATLSRX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATLSRX2H7L D GN Q QN RN SN VDD VSS
*.PININFO D:I GN:I RN:I SN:I Q:O QN:O VDD:B VSS:B
XI6 G VDD VSS GB / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI3 GN VDD VSS G / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI2 net0102 VDD VSS netqn / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI4 netqn VDD VSS QN / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI8 net0102 VDD VSS Q / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI1 SN VDD VSS S / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
MNM3 net0102 GB net41 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net0102 S VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM1 net47 D net44 VSS nm1p2_lvt_lp W=240n L=60n m=1
MNM2 net41 netqn net44 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM4 net44 RN VSS VSS nm1p2_lvt_lp W=240n L=60n m=1
XI7 G GB net47 net0102 VDD VSS / TG pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
MPM6 net053 netqn net059 VDD pm1p2_lvt_lp W=280n L=60n m=1
MPM4 net059 S VDD VDD pm1p2_lvt_lp W=340n L=60n m=1
MPM3 net47 D net059 VDD pm1p2_lvt_lp W=340n L=60n m=1
MPM0 net0102 RN net059 VDD pm1p2_lvt_lp W=200n L=60n m=1
MPM5 net0102 G net053 VDD pm1p2_lvt_lp W=280n L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATLSX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATLSX0P5H7L D GN Q QN SN VDD VSS
*.PININFO D:I GN:I SN:I Q:O QN:O VDD:B VSS:B
MNM1 net44 D VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM2 netq S VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM0 netq GB net38 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net38 netqn VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM4 net063 S VDD VDD pm1p2_lvt_lp W=320n L=60n m=1
MPM3 net44 D net063 VDD pm1p2_lvt_lp W=320n L=60n m=1
MPM2 net066 S VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM1 net057 netqn net066 VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM0 netq G net057 VDD pm1p2_lvt_lp W=150n L=60n m=1
XI0 netq VDD VSS Q / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI2 netq VDD VSS netqn / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI1 netqn VDD VSS QN / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI3 GN VDD VSS G / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI4 G VDD VSS GB / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI5 SN VDD VSS S / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI7 G GB net44 netq VDD VSS / TG pl=6E-08 pw=3.2E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATLSX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATLSX1H7L D GN Q QN SN VDD VSS
*.PININFO D:I GN:I SN:I Q:O QN:O VDD:B VSS:B
MNM1 net44 D VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM2 netq S VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM0 netq GB net38 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net38 netqn VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM4 net063 S VDD VDD pm1p2_lvt_lp W=320n L=60n m=1
MPM3 net44 D net063 VDD pm1p2_lvt_lp W=320n L=60n m=1
MPM2 net066 S VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM1 net057 netqn net066 VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM0 netq G net057 VDD pm1p2_lvt_lp W=150n L=60n m=1
XI0 netq VDD VSS Q / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI2 netq VDD VSS netqn / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI1 netqn VDD VSS QN / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI3 GN VDD VSS G / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI4 G VDD VSS GB / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI5 SN VDD VSS S / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI7 G GB net44 netq VDD VSS / TG pl=6E-08 pw=3.2E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATLSX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATLSX2H7L D GN Q QN SN VDD VSS
*.PININFO D:I GN:I SN:I Q:O QN:O VDD:B VSS:B
MNM1 net44 D VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM2 netq S VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM0 netq GB net38 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net38 netqn VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM4 net063 S VDD VDD pm1p2_lvt_lp W=320n L=60n m=1
MPM3 net44 D net063 VDD pm1p2_lvt_lp W=320n L=60n m=1
MPM2 net066 S VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM1 net057 netqn net066 VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM0 netq G net057 VDD pm1p2_lvt_lp W=150n L=60n m=1
XI0 netq VDD VSS Q / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI2 netq VDD VSS netqn / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI1 netqn VDD VSS QN / INV pl=6E-08 pw=4E-07 nl=6E-08 nw=2.8E-07
XI3 GN VDD VSS G / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI4 G VDD VSS GB / INV pl=6E-08 pw=3.4E-07 nl=6E-08 nw=2.4E-07
XI5 SN VDD VSS S / INV pl=6E-08 pw=2.8E-07 nl=6E-08 nw=2E-07
XI7 G GB net44 netq VDD VSS / TG pl=6E-08 pw=3.2E-07 nl=6E-08 nw=2E-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATLX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATLX0P5H7L D GN Q QN VDD VSS
*.PININFO D:I GN:I Q:O QN:O VDD:B VSS:B
XXI15 net9 GPN GP VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI6 D GP GPN VDD VSS net25 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI14 net9 VDD VSS QN / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XXI13 GP VDD VSS GPN / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net25 VDD VSS Q / INV pl=60n pw=280n nl=60n nw=200n
XXI4 GN VDD VSS GP / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATLX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATLX1H7L D GN Q QN VDD VSS
*.PININFO D:I GN:I Q:O QN:O VDD:B VSS:B
XXI15 net9 GPN GP VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI6 D GP GPN VDD VSS net25 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI7 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net25 VDD VSS Q / INV pl=60n pw=340n nl=60n nw=240n
XI0 net9 VDD VSS QN / INV pl=60n pw=340n nl=60n nw=240n
XXI13 GP VDD VSS GPN / INV pl=60n pw=280n nl=60n nw=200n
XXI4 GN VDD VSS GP / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATLX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATLX2H7L D GN Q QN VDD VSS
*.PININFO D:I GN:I Q:O QN:O VDD:B VSS:B
XXI6 D GP GPN VDD VSS net25 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI15 net9 GPN GP VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI7 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XXI4 GN VDD VSS GP / INV pl=60n pw=280n nl=60n nw=200n
XI0 net9 VDD VSS QN / INV pl=60n pw=400n nl=60n nw=280n
XXI13 GP VDD VSS GPN / INV pl=60n pw=280n nl=60n nw=200n
XI1 net25 VDD VSS Q / INV pl=60n pw=400n nl=60n nw=280n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATLX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATLX3H7L D GN Q QN VDD VSS
*.PININFO D:I GN:I Q:O QN:O VDD:B VSS:B
XXI15 net9 GPN GP VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI6 D GP GPN VDD VSS net25 / TSINV pl=60n pw=340n nl=60n nw=240n
XI0 net9 VDD VSS QN / INV pl=60n pw=600n nl=60n nw=420n
XI1 net25 VDD VSS Q / INV pl=60n pw=600n nl=60n nw=420n
XXI13 GP VDD VSS GPN / INV pl=60n pw=340n nl=60n nw=240n
XXI7 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XXI4 GN VDD VSS GP / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    LATLX4H7L
* View Name:    schematic
************************************************************************

.SUBCKT LATLX4H7L D GN Q QN VDD VSS
*.PININFO D:I GN:I Q:O QN:O VDD:B VSS:B
XXI6 D GP GPN VDD VSS net25 / TSINV pl=60n pw=340n nl=60n nw=240n
XXI15 net9 GPN GP VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI7 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XXI4 GN VDD VSS GP / INV pl=60n pw=280n nl=60n nw=200n
XI0 net9 VDD VSS QN / INV pl=60n pw=800n nl=60n nw=560n
XXI13 GP VDD VSS GPN / INV pl=60n pw=340n nl=60n nw=240n
XI2 net25 VDD VSS Q / INV pl=60n pw=800n nl=60n nw=560n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MDFFQX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT MDFFQX0P5H7L CK D0 D1 Q S0 VDD VSS
*.PININFO CK:I D0:I D1:I S0:I Q:O VDD:B VSS:B
XXI18 net32 net24 net030 net33 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
XXI14 net46 net24 net32 VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI17 D1 S0 net057 VDD VSS net030 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI19 D0 net057 S0 VDD VSS net030 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI9 net46 net24 net32 VDD VSS net25 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI15 net9 net32 net24 VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI20 S0 VDD VSS net057 / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=280n nl=60n nw=200n
XXI13 net32 VDD VSS net24 / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net25 VDD VSS Q / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XXI4 CK VDD VSS net32 / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MDFFQX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT MDFFQX1H7L CK D0 D1 Q S0 VDD VSS
*.PININFO CK:I D0:I D1:I S0:I Q:O VDD:B VSS:B
XXI18 net32 net24 net034 net33 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
XXI14 net46 net24 net32 VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI19 D1 S0 net057 VDD VSS net034 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI20 D0 net057 S0 VDD VSS net034 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI9 net46 net24 net32 VDD VSS net25 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI15 net9 net32 net24 VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI21 S0 VDD VSS net057 / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=280n nl=60n nw=200n
XXI13 net32 VDD VSS net24 / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net25 VDD VSS Q / INV pl=60n pw=340n nl=60n nw=240n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=300n nl=60n nw=220n
XXI4 CK VDD VSS net32 / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MDFFQX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT MDFFQX2H7L CK D0 D1 Q S0 VDD VSS
*.PININFO CK:I D0:I D1:I S0:I Q:O VDD:B VSS:B
XXI18 net32 net24 net034 net33 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
XXI14 net46 net24 net32 VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI19 D1 S0 net055 VDD VSS net034 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI20 D0 net055 S0 VDD VSS net034 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI9 net46 net24 net32 VDD VSS net25 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI15 net9 net32 net24 VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI21 S0 VDD VSS net055 / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=280n nl=60n nw=200n
XXI13 net32 VDD VSS net24 / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net25 VDD VSS Q / INV pl=60n pw=400n nl=60n nw=280n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=340n nl=60n nw=240n
XXI4 CK VDD VSS net32 / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MSDFFQX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT MSDFFQX0P5H7L CK D0 D1 Q S0 SE SI VDD VSS
*.PININFO CK:I D0:I D1:I S0:I SE:I SI:I Q:O VDD:B VSS:B
XXI21 c cn net46 net25 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
XXI20 SEN SE net034 net046 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
XXI14 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI24 D1 S0 S0N VDD VSS net034 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI25 D0 S0N S0 VDD VSS net034 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI22 SI SE SEN VDD VSS net046 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI19 net046 cn c VDD VSS net33 / TSINV pl=60n pw=300n nl=60n nw=220n
XXI15 net9 cn c VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI26 S0 VDD VSS S0N / INV pl=60n pw=280n nl=60n nw=200n
XXI23 SE VDD VSS SEN / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=280n nl=60n nw=200n
XXI13 cn VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net25 VDD VSS Q / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XXI4 CK VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MSDFFQX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT MSDFFQX1H7L CK D0 D1 Q S0 SE SI VDD VSS
*.PININFO CK:I D0:I D1:I S0:I SE:I SI:I Q:O VDD:B VSS:B
XXI21 c cn net46 net25 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
XXI20 SEN SE net034 net046 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
XXI14 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI24 D1 S0 S0N VDD VSS net034 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI25 D0 S0N S0 VDD VSS net034 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI22 SI SE SEN VDD VSS net046 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI19 net046 cn c VDD VSS net33 / TSINV pl=60n pw=300n nl=60n nw=220n
XXI15 net9 cn c VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI26 S0 VDD VSS S0N / INV pl=60n pw=280n nl=60n nw=200n
XXI23 SE VDD VSS SEN / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=300n nl=60n nw=220n
XXI13 cn VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net25 VDD VSS Q / INV pl=60n pw=340n nl=60n nw=240n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XXI4 CK VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MSDFFQX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT MSDFFQX2H7L CK D0 D1 Q S0 SE SI VDD VSS
*.PININFO CK:I D0:I D1:I S0:I SE:I SI:I Q:O VDD:B VSS:B
XXI20 SEN SE net034 net046 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
XXI21 c cn net46 net25 VDD VSS / TG pl=60n pw=340n nl=60n nw=240n
XXI15 net9 cn c VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI19 net046 cn c VDD VSS net33 / TSINV pl=60n pw=300n nl=60n nw=220n
XXI22 SI SE SEN VDD VSS net046 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI25 D0 S0N S0 VDD VSS net034 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI24 D1 S0 S0N VDD VSS net034 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI14 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI4 CK VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net25 VDD VSS Q / INV pl=60n pw=400n nl=60n nw=280n
XXI13 cn VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=340n nl=60n nw=240n
XXI23 SE VDD VSS SEN / INV pl=60n pw=280n nl=60n nw=200n
XXI26 S0 VDD VSS S0N / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MSDFFQX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT MSDFFQX3H7L CK D0 D1 Q S0 SE SI VDD VSS
*.PININFO CK:I D0:I D1:I S0:I SE:I SI:I Q:O VDD:B VSS:B
XXI22 SI SE SEN VDD VSS net046 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI15 net9 cn c VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI14 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI25 D0 S0N S0 VDD VSS net034 / TSINV pl=60n pw=310n nl=60n nw=220n
XXI19 net046 cn c VDD VSS net33 / TSINV pl=60n pw=320n nl=60n nw=230n
XXI24 D1 S0 S0N VDD VSS net034 / TSINV pl=60n pw=310n nl=60n nw=220n
XXI20 SEN SE net034 net046 VDD VSS / TG pl=60n pw=310n nl=60n nw=220n
XXI21 c cn net46 net25 VDD VSS / TG pl=60n pw=350n nl=60n nw=250n
XXI4 CK VDD VSS cn / INV pl=60n pw=295n nl=60n nw=210n
XXI13 cn VDD VSS c / INV pl=60n pw=295n nl=60n nw=210n
XXI23 SE VDD VSS SEN / INV pl=60n pw=310n nl=60n nw=220n
XXI26 S0 VDD VSS S0N / INV pl=60n pw=310n nl=60n nw=220n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=350n nl=60n nw=250n
XXI12 net25 VDD VSS Q / INV pl=60n pw=600n nl=60n nw=420n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUX2X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUX2X0P5H7L A B S0 VDD VSS Y
*.PININFO A:I B:I S0:I Y:O VDD:B VSS:B
XXI2 net19 VDD VSS Y / INV pl=60n pw=190n nl=60n nw=150n
XXI0 S0 VDD VSS S0N / INV pl=60n pw=190n nl=60n nw=150n
XXI5 B S0 S0N VDD VSS net19 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI3 A S0N S0 VDD VSS net19 / TSINV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUX2X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUX2X0P7H7L A B S0 VDD VSS Y
*.PININFO A:I B:I S0:I Y:O VDD:B VSS:B
XXI0 S0 VDD VSS S0N / INV pl=60n pw=190n nl=60n nw=150n
XXI2 net19 VDD VSS Y / INV pl=60n pw=222n nl=60n nw=174n
XXI3 A S0N S0 VDD VSS net19 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI5 B S0 S0N VDD VSS net19 / TSINV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUX2X12H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUX2X12H7L A B S0 VDD VSS Y
*.PININFO A:I B:I S0:I Y:O VDD:B VSS:B
XXI9 B VDD VSS BN / INV pl=60n pw=930n nl=60n nw=750n
XXI7 A VDD VSS AN / INV pl=60n pw=930n nl=60n nw=750n
XXI0 S0 VDD VSS S0N / INV pl=60n pw=380n nl=60n nw=300n
XXI2 net19 VDD VSS Y / INV pl=60n pw=2.28u nl=60n nw=1.8u
XXI8 S0 S0N BN net19 VDD VSS / TG pl=60n pw=930n nl=60n nw=750n
XXI6 S0N S0 AN net19 VDD VSS / TG pl=60n pw=930n nl=60n nw=750n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUX2X16H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUX2X16H7L A B S0 VDD VSS Y
*.PININFO A:I B:I S0:I Y:O VDD:B VSS:B
XXI9 B VDD VSS BN / INV pl=60n pw=1.24u nl=60n nw=1u
XXI7 A VDD VSS AN / INV pl=60n pw=1.24u nl=60n nw=1u
XXI0 S0 VDD VSS S0N / INV pl=60n pw=380n nl=60n nw=300n
XXI2 net19 VDD VSS Y / INV pl=60n pw=3.04u nl=60n nw=2.4u
XXI8 S0 S0N BN net19 VDD VSS / TG pl=60n pw=1.24u nl=60n nw=1u
XXI6 S0N S0 AN net19 VDD VSS / TG pl=60n pw=1.24u nl=60n nw=1u
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUX2X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUX2X1H7L A B S0 VDD VSS Y
*.PININFO A:I B:I S0:I Y:O VDD:B VSS:B
XXI0 S0 VDD VSS S0N / INV pl=60n pw=190n nl=60n nw=150n
XXI2 net19 VDD VSS Y / INV pl=60n pw=270n nl=60n nw=210n
XXI3 A S0N S0 VDD VSS net19 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI5 B S0 S0N VDD VSS net19 / TSINV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUX2X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUX2X1P4H7L A B S0 VDD VSS Y
*.PININFO A:I B:I S0:I Y:O VDD:B VSS:B
XXI0 S0 VDD VSS S0N / INV pl=60n pw=190n nl=60n nw=150n
XXI2 net19 VDD VSS Y / INV pl=60n pw=314n nl=60n nw=246n
XXI3 A S0N S0 VDD VSS net19 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI5 B S0 S0N VDD VSS net19 / TSINV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUX2X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUX2X2H7L A B S0 VDD VSS Y
*.PININFO A:I B:I S0:I Y:O VDD:B VSS:B
XXI9 B VDD VSS BN / INV pl=60n pw=190n nl=60n nw=150n
XXI7 A VDD VSS AN / INV pl=60n pw=190n nl=60n nw=150n
XXI0 S0 VDD VSS S0N / INV pl=60n pw=190n nl=60n nw=150n
XXI2 net19 VDD VSS Y / INV pl=60n pw=380n nl=60n nw=300n
XXI8 S0 S0N BN net19 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI6 S0N S0 AN net19 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUX2X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUX2X3H7L A B S0 VDD VSS Y
*.PININFO A:I B:I S0:I Y:O VDD:B VSS:B
XXI2 net19 VDD VSS Y / INV pl=60n pw=570n nl=60n nw=450n
XXI0 S0 VDD VSS S0N / INV pl=60n pw=200n nl=60n nw=160n
XXI7 A VDD VSS AN / INV pl=60n pw=250n nl=60n nw=200n
XXI9 B VDD VSS BN / INV pl=60n pw=250n nl=60n nw=200n
XXI6 S0N S0 AN net19 VDD VSS / TG pl=60n pw=250n nl=60n nw=200n
XXI8 S0 S0N BN net19 VDD VSS / TG pl=60n pw=250n nl=60n nw=200n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUX2X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUX2X4H7L A B S0 VDD VSS Y
*.PININFO A:I B:I S0:I Y:O VDD:B VSS:B
XXI9 B VDD VSS BN / INV pl=60n pw=310n nl=60n nw=250n
XXI7 A VDD VSS AN / INV pl=60n pw=310n nl=60n nw=250n
XXI0 S0 VDD VSS S0N / INV pl=60n pw=210n nl=60n nw=170n
XXI2 net19 VDD VSS Y / INV pl=60n pw=760n nl=60n nw=600n
XXI8 S0 S0N BN net19 VDD VSS / TG pl=60n pw=310n nl=60n nw=250n
XXI6 S0N S0 AN net19 VDD VSS / TG pl=60n pw=310n nl=60n nw=250n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUX2X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUX2X6H7L A B S0 VDD VSS Y
*.PININFO A:I B:I S0:I Y:O VDD:B VSS:B
XXI9 B VDD VSS BN / INV pl=60n pw=380n nl=60n nw=300n
XXI7 A VDD VSS AN / INV pl=60n pw=380n nl=60n nw=300n
XXI0 S0 VDD VSS S0N / INV pl=60n pw=250n nl=60n nw=200n
XXI2 net19 VDD VSS Y / INV pl=60n pw=1140n nl=60n nw=900n
XXI8 S0 S0N BN net19 VDD VSS / TG pl=60n pw=380n nl=60n nw=300n
XXI6 S0N S0 AN net19 VDD VSS / TG pl=60n pw=380n nl=60n nw=300n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUX2X8H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUX2X8H7L A B S0 VDD VSS Y
*.PININFO A:I B:I S0:I Y:O VDD:B VSS:B
XXI9 B VDD VSS BN / INV pl=60n pw=620n nl=60n nw=500n
XXI7 A VDD VSS AN / INV pl=60n pw=620n nl=60n nw=500n
XXI0 S0 VDD VSS S0N / INV pl=60n pw=380n nl=60n nw=300n
XXI2 net19 VDD VSS Y / INV pl=60n pw=1520n nl=60n nw=1200n
XXI8 S0 S0N BN net19 VDD VSS / TG pl=60n pw=620n nl=60n nw=500n
XXI6 S0N S0 AN net19 VDD VSS / TG pl=60n pw=620n nl=60n nw=500n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUX4X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUX4X0P5H7L A B C D S0 S1 VDD VSS Y
*.PININFO A:I B:I C:I D:I S0:I S1:I Y:O VDD:B VSS:B
XXI9 S1 VDD VSS S1N / INV pl=60n pw=190n nl=60n nw=150n
XXI8 S0 VDD VSS S0N / INV pl=60n pw=190n nl=60n nw=150n
XXI1 net9 VDD VSS Y / INV pl=60n pw=190n nl=60n nw=150n
XXI10 S1N S1 net25 net9 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI11 S1 S1N net17 net9 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI7 D S0 S0N VDD VSS net17 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI6 C S0N S0 VDD VSS net17 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI5 B S0 S0N VDD VSS net25 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI4 A S0N S0 VDD VSS net25 / TSINV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUX4X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUX4X0P7H7L A B C D S0 S1 VDD VSS Y
*.PININFO A:I B:I C:I D:I S0:I S1:I Y:O VDD:B VSS:B
XXI9 S1 VDD VSS S1N / INV pl=60n pw=190n nl=60n nw=150n
XXI8 S0 VDD VSS S0N / INV pl=60n pw=190n nl=60n nw=150n
XXI1 net9 VDD VSS Y / INV pl=60n pw=222n nl=60n nw=174n
XXI10 S1N S1 net25 net9 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI11 S1 S1N net17 net9 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI7 D S0 S0N VDD VSS net17 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI6 C S0N S0 VDD VSS net17 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI5 B S0 S0N VDD VSS net25 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI4 A S0N S0 VDD VSS net25 / TSINV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUX4X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUX4X1H7L A B C D S0 S1 VDD VSS Y
*.PININFO A:I B:I C:I D:I S0:I S1:I Y:O VDD:B VSS:B
XXI9 S1 VDD VSS S1N / INV pl=60n pw=190n nl=60n nw=150n
XXI8 S0 VDD VSS S0N / INV pl=60n pw=190n nl=60n nw=150n
XXI1 net9 VDD VSS Y / INV pl=60n pw=270n nl=60n nw=210n
XXI10 S1N S1 net25 net9 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI11 S1 S1N net17 net9 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI7 D S0 S0N VDD VSS net17 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI6 C S0N S0 VDD VSS net17 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI5 B S0 S0N VDD VSS net25 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI4 A S0N S0 VDD VSS net25 / TSINV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUX4X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUX4X1P4H7L A B C D S0 S1 VDD VSS Y
*.PININFO A:I B:I C:I D:I S0:I S1:I Y:O VDD:B VSS:B
XXI9 S1 VDD VSS S1N / INV pl=60n pw=190n nl=60n nw=150n
XXI8 S0 VDD VSS S0N / INV pl=60n pw=190n nl=60n nw=150n
XXI1 net9 VDD VSS Y / INV pl=60n pw=314n nl=60n nw=246n
XXI10 S1N S1 net25 net9 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI11 S1 S1N net17 net9 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI7 D S0 S0N VDD VSS net17 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI6 C S0N S0 VDD VSS net17 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI5 B S0 S0N VDD VSS net25 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI4 A S0N S0 VDD VSS net25 / TSINV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUX4X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUX4X2H7L A B C D S0 S1 VDD VSS Y
*.PININFO A:I B:I C:I D:I S0:I S1:I Y:O VDD:B VSS:B
XXI9 S1 VDD VSS S1N / INV pl=60n pw=190n nl=60n nw=150n
XXI8 S0 VDD VSS S0N / INV pl=60n pw=190n nl=60n nw=150n
XXI1 net9 VDD VSS Y / INV pl=60n pw=380n nl=60n nw=300n
XXI10 S1N S1 net25 net9 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI11 S1 S1N net17 net9 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI7 D S0 S0N VDD VSS net17 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI6 C S0N S0 VDD VSS net17 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI5 B S0 S0N VDD VSS net25 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI4 A S0N S0 VDD VSS net25 / TSINV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUX4X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUX4X3H7L A B C D S0 S1 VDD VSS Y
*.PININFO A:I B:I C:I D:I S0:I S1:I Y:O VDD:B VSS:B
XXI1 net9 VDD VSS Y / INV pl=60n pw=570n nl=60n nw=450n
XXI8 S0 VDD VSS S0N / INV pl=60n pw=250n nl=60n nw=200n
XXI9 S1 VDD VSS S1N / INV pl=60n pw=195n nl=60n nw=160n
XXI11 S1 S1N net17 net9 VDD VSS / TG pl=60n pw=250n nl=60n nw=200n
XXI10 S1N S1 net25 net9 VDD VSS / TG pl=60n pw=250n nl=60n nw=200n
XXI4 A S0N S0 VDD VSS net25 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI5 B S0 S0N VDD VSS net25 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI6 C S0N S0 VDD VSS net17 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI7 D S0 S0N VDD VSS net17 / TSINV pl=60n pw=250n nl=60n nw=200n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUX4X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUX4X4H7L A B C D S0 S1 VDD VSS Y
*.PININFO A:I B:I C:I D:I S0:I S1:I Y:O VDD:B VSS:B
XXI1 net9 VDD VSS Y / INV pl=60n pw=760n nl=60n nw=600n
XXI8 S0 VDD VSS S0N / INV pl=60n pw=310n nl=60n nw=250n
XXI9 S1 VDD VSS S1N / INV pl=60n pw=200n nl=60n nw=170n
XXI11 S1 S1N net17 net9 VDD VSS / TG pl=60n pw=310n nl=60n nw=250n
XXI10 S1N S1 net25 net9 VDD VSS / TG pl=60n pw=310n nl=60n nw=250n
XXI4 A S0N S0 VDD VSS net25 / TSINV pl=60n pw=310n nl=60n nw=250n
XXI5 B S0 S0N VDD VSS net25 / TSINV pl=60n pw=310n nl=60n nw=250n
XXI6 C S0N S0 VDD VSS net17 / TSINV pl=60n pw=310n nl=60n nw=250n
XXI7 D S0 S0N VDD VSS net17 / TSINV pl=60n pw=310n nl=60n nw=250n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUX4X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUX4X6H7L A B C D S0 S1 VDD VSS Y
*.PININFO A:I B:I C:I D:I S0:I S1:I Y:O VDD:B VSS:B
XXI1 net9 VDD VSS Y / INV pl=60n pw=1.14u nl=60n nw=0.9u
XXI8 S0 VDD VSS S0N / INV pl=60n pw=380n nl=60n nw=300n
XXI9 S1 VDD VSS S1N / INV pl=60n pw=250n nl=60n nw=200n
XXI11 S1 S1N net17 net9 VDD VSS / TG pl=60n pw=310n nl=60n nw=250n
XXI10 S1N S1 net25 net9 VDD VSS / TG pl=60n pw=310n nl=60n nw=250n
XXI4 A S0N S0 VDD VSS net25 / TSINV pl=60n pw=380n nl=60n nw=300n
XXI5 B S0 S0N VDD VSS net25 / TSINV pl=60n pw=380n nl=60n nw=300n
XXI6 C S0N S0 VDD VSS net17 / TSINV pl=60n pw=380n nl=60n nw=300n
XXI7 D S0 S0N VDD VSS net17 / TSINV pl=60n pw=380n nl=60n nw=300n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUXI2X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUXI2X0P5H7L A B S0 VDD VSS Y
*.PININFO A:I B:I S0:I Y:O VDD:B VSS:B
XXI9 A VDD VSS net030 / INV pl=60n pw=190n nl=60n nw=150n
XXI10 B VDD VSS net028 / INV pl=60n pw=190n nl=60n nw=150n
XXI0 S0 VDD VSS S0N / INV pl=60n pw=190n nl=60n nw=150n
XXI8 S0 S0N net028 Y VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI7 S0N S0 net030 Y VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUXI2X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUXI2X0P7H7L A B S0 VDD VSS Y
*.PININFO A:I B:I S0:I Y:O VDD:B VSS:B
XXI9 A VDD VSS net030 / INV pl=60n pw=222n nl=60n nw=174n
XXI10 B VDD VSS net028 / INV pl=60n pw=222n nl=60n nw=174n
XXI0 S0 VDD VSS S0N / INV pl=60n pw=190n nl=60n nw=150n
XXI8 S0 S0N net028 Y VDD VSS / TG pl=60n pw=222n nl=60n nw=174n
XXI7 S0N S0 net030 Y VDD VSS / TG pl=60n pw=222n nl=60n nw=174n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUXI2X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUXI2X1H7L A B S0 VDD VSS Y
*.PININFO A:I B:I S0:I Y:O VDD:B VSS:B
XXI9 A VDD VSS net030 / INV pl=60n pw=270n nl=60n nw=210n
XXI10 B VDD VSS net028 / INV pl=60n pw=270n nl=60n nw=210n
XXI0 S0 VDD VSS S0N / INV pl=60n pw=190n nl=60n nw=150n
XXI8 S0 S0N net028 Y VDD VSS / TG pl=60n pw=270n nl=60n nw=210n
XXI7 S0N S0 net030 Y VDD VSS / TG pl=60n pw=270n nl=60n nw=210n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUXI2X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUXI2X1P4H7L A B S0 VDD VSS Y
*.PININFO A:I B:I S0:I Y:O VDD:B VSS:B
XXI9 A VDD VSS net030 / INV pl=60n pw=314n nl=60n nw=246n
XXI10 B VDD VSS net028 / INV pl=60n pw=314n nl=60n nw=246n
XXI0 S0 VDD VSS S0N / INV pl=60n pw=190n nl=60n nw=150n
XXI8 S0 S0N net028 Y VDD VSS / TG pl=60n pw=314n nl=60n nw=246n
XXI7 S0N S0 net030 Y VDD VSS / TG pl=60n pw=314n nl=60n nw=246n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUXI2X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUXI2X2H7L A B S0 VDD VSS Y
*.PININFO A:I B:I S0:I Y:O VDD:B VSS:B
XXI7 S0N S0 net030 Y VDD VSS / TG pl=60n pw=380n nl=60n nw=300n
XXI8 S0 S0N net028 Y VDD VSS / TG pl=60n pw=380n nl=60n nw=300n
XXI0 S0 VDD VSS S0N / INV pl=60n pw=190n nl=60n nw=150n
XXI10 B VDD VSS net028 / INV pl=60n pw=380n nl=60n nw=300n
XXI9 A VDD VSS net030 / INV pl=60n pw=380n nl=60n nw=300n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUXI2X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUXI2X3H7L A B S0 VDD VSS Y
*.PININFO A:I B:I S0:I Y:O VDD:B VSS:B
XXI8 S0 S0N net028 Y VDD VSS / TG pl=60n pw=510n nl=60n nw=435n
XXI7 S0N S0 net030 Y VDD VSS / TG pl=60n pw=510n nl=60n nw=435n
XXI0 S0 VDD VSS S0N / INV pl=60n pw=250n nl=60n nw=200n
XXI9 A VDD VSS net030 / INV pl=60n pw=570n nl=60n nw=450n
XXI10 B VDD VSS net028 / INV pl=60n pw=570n nl=60n nw=450n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    MUXI2X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT MUXI2X4H7L A B S0 VDD VSS Y
*.PININFO A:I B:I S0:I Y:O VDD:B VSS:B
XXI8 S0 S0N net028 Y VDD VSS / TG pl=60n pw=640n nl=60n nw=570n
XXI7 S0N S0 net030 Y VDD VSS / TG pl=60n pw=640n nl=60n nw=570n
XXI0 S0 VDD VSS S0N / INV pl=60n pw=310n nl=60n nw=250n
XXI9 A VDD VSS net030 / INV pl=60n pw=760n nl=60n nw=600n
XXI10 B VDD VSS net028 / INV pl=60n pw=760n nl=60n nw=600n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND2BX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2BX0P5H7L AN B VDD VSS Y
*.PININFO AN:I B:I Y:O VDD:B VSS:B
MMN0 Y B net6 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 net6 net14 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP1 Y net14 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 AN VDD VSS net14 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND2BX0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2BX0P7H7L AN B VDD VSS Y
*.PININFO AN:I B:I Y:O VDD:B VSS:B
MMN0 Y B net6 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN1 net6 net036 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMP1 Y net036 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
XXI3 AN VDD VSS net036 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND2BX12H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2BX12H7L AN B VDD VSS Y
*.PININFO AN:I B:I Y:O VDD:B VSS:B
MMM4 net16 AN VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMM1 Y B VDD VDD pm1p2_lvt_lp W=2.28u L=60n m=1
MMM0 Y net16 VDD VDD pm1p2_lvt_lp W=2.28u L=60n m=1
MMM5 net16 AN VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMM2 net20 net16 VSS VSS nm1p2_lvt_lp W=1.8u L=60n m=1
MMM3 Y B net20 VSS nm1p2_lvt_lp W=1.8u L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND2BX16H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2BX16H7L AN B VDD VSS Y
*.PININFO AN:I B:I Y:O VDD:B VSS:B
MMM5 net16 AN VSS VSS nm1p2_lvt_lp W=2.4u L=60n m=1
MMM2 net20 net16 VSS VSS nm1p2_lvt_lp W=2.4u L=60n m=1
MMM3 Y B net20 VSS nm1p2_lvt_lp W=2.4u L=60n m=1
MMM4 net16 AN VDD VDD pm1p2_lvt_lp W=3.04u L=60n m=1
MMM1 Y B VDD VDD pm1p2_lvt_lp W=3.04u L=60n m=1
MMM0 Y net16 VDD VDD pm1p2_lvt_lp W=3.04u L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND2BX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2BX1H7L AN B VDD VSS Y
*.PININFO AN:I B:I Y:O VDD:B VSS:B
MMN0 Y B net6 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN1 net6 net036 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMP1 Y net036 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
XXI3 AN VDD VSS net036 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND2BX1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2BX1P4H7L AN B VDD VSS Y
*.PININFO AN:I B:I Y:O VDD:B VSS:B
MMN0 Y B net6 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN1 net6 net036 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMP1 Y net036 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
XXI3 AN VDD VSS net036 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND2BX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2BX2H7L AN B VDD VSS Y
*.PININFO AN:I B:I Y:O VDD:B VSS:B
MMN0 Y B net6 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN1 net6 net14 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP1 Y net14 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
XXI3 AN VDD VSS net14 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND2BX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2BX3H7L AN B VDD VSS Y
*.PININFO AN:I B:I Y:O VDD:B VSS:B
MMN0 Y B net6 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN1 net6 net036 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMP1 Y net036 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
XXI3 AN VDD VSS net036 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND2BX4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2BX4H7L AN B VDD VSS Y
*.PININFO AN:I B:I Y:O VDD:B VSS:B
MMN0 Y B net6 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN1 net6 net14 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMP1 Y net14 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
XXI3 AN VDD VSS net14 / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND2BX6H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2BX6H7L AN B VDD VSS Y
*.PININFO AN:I B:I Y:O VDD:B VSS:B
MMM4 net16 AN VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMM1 Y B VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMM0 Y net16 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMM5 net16 AN VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMM2 net20 net16 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMM3 Y B net20 VSS nm1p2_lvt_lp W=900n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND2BX8H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2BX8H7L AN B VDD VSS Y
*.PININFO AN:I B:I Y:O VDD:B VSS:B
MMM4 net16 AN VDD VDD pm1p2_lvt_lp W=620n L=60n m=1
MMM1 Y B VDD VDD pm1p2_lvt_lp W=1.52u L=60n m=1
MMM0 Y net16 VDD VDD pm1p2_lvt_lp W=1.52u L=60n m=1
MMM5 net16 AN VSS VSS nm1p2_lvt_lp W=500n L=60n m=1
MMM2 net20 net16 VSS VSS nm1p2_lvt_lp W=1.2u L=60n m=1
MMM3 Y B net20 VSS nm1p2_lvt_lp W=1.2u L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND2X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2X0P5H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net6 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 net6 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP0 Y A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND2X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2X0P7H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net6 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN1 net6 A VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP0 Y A VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND2X12H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2X12H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMM3 Y B net12 VSS nm1p2_lvt_lp W=1.8u L=60n m=1
MMM2 net12 A VSS VSS nm1p2_lvt_lp W=1.8u L=60n m=1
MMM1 Y B VDD VDD pm1p2_lvt_lp W=2.28u L=60n m=1
MMM0 Y A VDD VDD pm1p2_lvt_lp W=2.28u L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND2X16H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2X16H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMM1 Y B VDD VDD pm1p2_lvt_lp W=3.04u L=60n m=1
MMM0 Y A VDD VDD pm1p2_lvt_lp W=3.04u L=60n m=1
MMM3 Y B net12 VSS nm1p2_lvt_lp W=2.4u L=60n m=1
MMM2 net12 A VSS VSS nm1p2_lvt_lp W=2.4u L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND2X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2X1H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net6 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN1 net6 A VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP0 Y A VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND2X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2X1P4H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net6 VSS nm1p2_lvt_lp W=246n L=60n m=1
MMN1 net6 A VSS VSS nm1p2_lvt_lp W=246n L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP0 Y A VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND2X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2X2H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net6 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN1 net6 A VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP0 Y A VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND2X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2X3H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net6 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN1 net6 A VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP0 Y A VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND2X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2X4H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net6 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN1 net6 A VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP0 Y A VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND2X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2X6H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMM3 Y B net12 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMM2 net12 A VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMM1 Y B VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMM0 Y A VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND2X8H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2X8H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMM1 Y B VDD VDD pm1p2_lvt_lp W=1.52u L=60n m=1
MMM0 Y A VDD VDD pm1p2_lvt_lp W=1.52u L=60n m=1
MMM3 Y B net12 VSS nm1p2_lvt_lp W=1.2u L=60n m=1
MMM2 net12 A VSS VSS nm1p2_lvt_lp W=1.2u L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3BBX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3BBX0P5H7L AN BN C VDD VSS Y
*.PININFO AN:I BN:I C:I Y:O VDD:B VSS:B
MMM2 net25 A2N net33 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM3 Y A1N net25 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM7 net33 C VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM5 A2N BN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM8 A1N AN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM1 Y C VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM0 Y A2N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM6 Y A1N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM4 A2N BN VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM9 A1N AN VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3BBX0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3BBX0P7H7L AN BN C VDD VSS Y
*.PININFO AN:I BN:I C:I Y:O VDD:B VSS:B
MMM2 net25 A2N net33 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMM3 Y A1N net25 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMM7 net33 C VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMM5 A2N BN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM8 A1N AN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM1 Y C VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMM0 Y A2N VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMM6 Y A1N VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMM4 A2N BN VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM9 A1N AN VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3BBX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3BBX1H7L AN BN C VDD VSS Y
*.PININFO AN:I BN:I C:I Y:O VDD:B VSS:B
MMM2 net25 A2N net33 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMM3 Y A1N net25 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMM7 net33 C VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMM5 A2N BN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM8 A1N AN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM1 Y C VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMM0 Y A2N VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMM6 Y A1N VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMM4 A2N BN VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM9 A1N AN VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3BBX1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3BBX1P4H7L AN BN C VDD VSS Y
*.PININFO AN:I BN:I C:I Y:O VDD:B VSS:B
MMM2 net25 A2N net33 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMM3 Y A1N net25 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMM7 net33 C VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMM5 A2N BN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM8 A1N AN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM1 Y C VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMM0 Y A2N VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMM6 Y A1N VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMM4 A2N BN VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM9 A1N AN VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3BBX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3BBX2H7L AN BN C VDD VSS Y
*.PININFO AN:I BN:I C:I Y:O VDD:B VSS:B
MMM2 net25 A2N net33 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM3 Y A1N net25 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM7 net33 C VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM5 A2N BN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM8 A1N AN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM1 Y C VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMM0 Y A2N VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMM6 Y A1N VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMM4 A2N BN VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMM9 A1N AN VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3BBX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3BBX3H7L AN BN C VDD VSS Y
*.PININFO AN:I BN:I C:I Y:O VDD:B VSS:B
MMM2 net25 A2N net33 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMM3 Y A1N net25 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMM7 net33 C VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMM5 A2N BN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM8 A1N AN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM1 Y C VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMM0 Y A2N VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMM6 Y A1N VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMM4 A2N BN VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM9 A1N AN VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3BBX4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3BBX4H7L AN BN C VDD VSS Y
*.PININFO AN:I BN:I C:I Y:O VDD:B VSS:B
MMM2 net25 A2N net33 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMM3 Y A1N net25 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMM7 net33 C VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMM5 A2N BN VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMM8 A1N AN VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMM1 Y C VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMM0 Y A2N VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMM6 Y A1N VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMM4 A2N BN VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMM9 A1N AN VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3BBX6H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3BBX6H7L AN BN C VDD VSS Y
*.PININFO AN:I BN:I C:I Y:O VDD:B VSS:B
MMM2 net25 A2N net33 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMM3 Y A1N net25 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMM7 net33 C VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMM5 A2N BN VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMM8 A1N AN VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMM1 Y C VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMM0 Y A2N VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMM6 Y A1N VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMM4 A2N BN VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMM9 A1N AN VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3BX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3BX0P5H7L AN B C VDD VSS Y
*.PININFO AN:I B:I C:I Y:O VDD:B VSS:B
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net7 net20 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 Y C net10 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP2 Y C VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP0 Y net20 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 AN VDD VSS net20 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3BX0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3BX0P7H7L AN B C VDD VSS Y
*.PININFO AN:I B:I C:I Y:O VDD:B VSS:B
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN4 net7 net20 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN0 Y C net10 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMP2 Y C VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP0 Y net20 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
XXI3 AN VDD VSS net20 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3BX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3BX1H7L AN B C VDD VSS Y
*.PININFO AN:I B:I C:I Y:O VDD:B VSS:B
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN4 net7 net20 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN0 Y C net10 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMP2 Y C VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP0 Y net20 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
XXI3 AN VDD VSS net20 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3BX1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3BX1P4H7L AN B C VDD VSS Y
*.PININFO AN:I B:I C:I Y:O VDD:B VSS:B
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN4 net7 net20 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN0 Y C net10 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMP2 Y C VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP0 Y net20 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
XXI3 AN VDD VSS net20 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3BX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3BX2H7L AN B C VDD VSS Y
*.PININFO AN:I B:I C:I Y:O VDD:B VSS:B
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN4 net7 net20 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN0 Y C net10 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP2 Y C VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP0 Y net20 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
XXI3 AN VDD VSS net20 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3BX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3BX3H7L AN B C VDD VSS Y
*.PININFO AN:I B:I C:I Y:O VDD:B VSS:B
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN4 net7 net20 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN0 Y C net10 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMP2 Y C VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP0 Y net20 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
XXI3 AN VDD VSS net20 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3BX4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3BX4H7L AN B C VDD VSS Y
*.PININFO AN:I B:I C:I Y:O VDD:B VSS:B
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN4 net7 net20 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN0 Y C net10 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMP2 Y C VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP0 Y net20 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
XXI3 AN VDD VSS net20 / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3BX6H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3BX6H7L AN B C VDD VSS Y
*.PININFO AN:I B:I C:I Y:O VDD:B VSS:B
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN4 net7 net20 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN0 Y C net10 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMP2 Y C VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP0 Y net20 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
XXI3 AN VDD VSS net20 / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3X0P5H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net7 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 Y C net10 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP2 Y C VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP0 Y A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3X0P7H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN4 net7 A VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN0 Y C net10 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMP2 Y C VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP0 Y A VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3X1H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN4 net7 A VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN0 Y C net10 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMP2 Y C VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP0 Y A VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3X1P4H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN4 net7 A VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN0 Y C net10 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMP2 Y C VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP0 Y A VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3X2H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN4 net7 A VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN0 Y C net10 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP2 Y C VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP0 Y A VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3X3H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN4 net7 A VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN0 Y C net10 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMP2 Y C VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP0 Y A VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3X4H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN4 net7 A VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN0 Y C net10 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMP2 Y C VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP0 Y A VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3X6H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN4 net7 A VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN0 Y C net10 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMP2 Y C VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP0 Y A VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND3X8H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3X8H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN3 net10 B net7 VSS nm1p2_lvt_lp W=1.2u L=60n m=1
MMN4 net7 A VSS VSS nm1p2_lvt_lp W=1.2u L=60n m=1
MMN0 Y C net10 VSS nm1p2_lvt_lp W=1.2u L=60n m=1
MMP2 Y C VDD VDD pm1p2_lvt_lp W=1.52u L=60n m=1
MMP1 Y B VDD VDD pm1p2_lvt_lp W=1.52u L=60n m=1
MMP0 Y A VDD VDD pm1p2_lvt_lp W=1.52u L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4BBX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4BBX0P5H7L AN BN C D VDD VSS Y
*.PININFO AN:I BN:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 net39 net32 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net32 net42 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP3 Y net42 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP0 Y net39 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI5 BN VDD VSS net39 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI6 AN VDD VSS net42 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4BBX0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4BBX0P7H7L AN BN C D VDD VSS Y
*.PININFO AN:I BN:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 net39 net32 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN5 net32 net42 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMP3 Y net42 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP0 Y net39 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
XXI5 BN VDD VSS net39 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI6 AN VDD VSS net42 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4BBX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4BBX1H7L AN BN C D VDD VSS Y
*.PININFO AN:I BN:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 net39 net32 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN5 net32 net42 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMP3 Y net42 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP0 Y net39 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
XXI5 BN VDD VSS net39 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI6 AN VDD VSS net42 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4BBX1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4BBX1P4H7L AN BN C D VDD VSS Y
*.PININFO AN:I BN:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 net39 net32 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN5 net32 net42 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMP3 Y net42 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP0 Y net39 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
XXI5 BN VDD VSS net39 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI6 AN VDD VSS net42 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4BBX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4BBX2H7L AN BN C D VDD VSS Y
*.PININFO AN:I BN:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 net39 net32 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN5 net32 net42 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP3 Y net42 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP0 Y net39 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
XXI5 BN VDD VSS net39 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI6 AN VDD VSS net42 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4BBX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4BBX3H7L AN BN C D VDD VSS Y
*.PININFO AN:I BN:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 net39 net32 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN5 net32 net42 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMP3 Y net42 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP0 Y net39 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
XXI5 BN VDD VSS net39 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI6 AN VDD VSS net42 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4BBX4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4BBX4H7L AN BN C D VDD VSS Y
*.PININFO AN:I BN:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 net39 net32 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN5 net32 net42 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMP3 Y net42 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP0 Y net39 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
XXI5 BN VDD VSS net39 / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
XXI6 AN VDD VSS net42 / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4BBX6H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4BBX6H7L AN BN C D VDD VSS Y
*.PININFO AN:I BN:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 net39 net32 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN5 net32 net42 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMP3 Y net42 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP0 Y net39 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
XXI5 BN VDD VSS net39 / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
XXI6 AN VDD VSS net42 / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4BX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4BX0P5H7L AN B C D VDD VSS Y
*.PININFO AN:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 B net28 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net28 net36 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP3 Y net36 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 AN VDD VSS net36 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4BX0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4BX0P7H7L AN B C D VDD VSS Y
*.PININFO AN:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 B net28 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN5 net28 net36 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMP3 Y net36 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
XXI3 AN VDD VSS net36 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4BX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4BX1H7L AN B C D VDD VSS Y
*.PININFO AN:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 B net28 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN5 net28 net36 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMP3 Y net36 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
XXI3 AN VDD VSS net36 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4BX1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4BX1P4H7L AN B C D VDD VSS Y
*.PININFO AN:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 B net28 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN5 net28 net36 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMP3 Y net36 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
XXI3 AN VDD VSS net36 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4BX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4BX2H7L AN B C D VDD VSS Y
*.PININFO AN:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 B net28 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN5 net28 net36 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP3 Y net36 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
XXI3 AN VDD VSS net36 / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4BX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4BX3H7L AN B C D VDD VSS Y
*.PININFO AN:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 B net28 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN5 net28 net36 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMP3 Y net36 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
XXI3 AN VDD VSS net36 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4BX4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4BX4H7L AN B C D VDD VSS Y
*.PININFO AN:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 B net28 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN5 net28 net36 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMP3 Y net36 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
XXI3 AN VDD VSS net36 / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4BX6H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4BX6H7L AN B C D VDD VSS Y
*.PININFO AN:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 B net28 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN5 net28 net36 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMP3 Y net36 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
XXI3 AN VDD VSS net36 / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4X0P5H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 B net25 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net25 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP3 Y A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4X0P7H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 B net25 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN5 net25 A VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMP3 Y A VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4X1H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 B net25 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN5 net25 A VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMP3 Y A VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4X1P4H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 B net25 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN5 net25 A VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMP3 Y A VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4X2H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 B net25 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN5 net25 A VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP3 Y A VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4X3H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 B net25 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN5 net25 A VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMP3 Y A VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4X4H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 B net25 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN5 net25 A VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMP3 Y A VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NAND4X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4X6H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 net7 B net25 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN5 net25 A VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN3 net10 C net7 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN0 Y D net10 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMP3 Y A VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP2 Y D VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP1 Y C VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR2BX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2BX0P5H7L AN B VDD VSS Z
*.PININFO AN:I B:I Z:O VDD:B VSS:B
MMN2 Z B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 Z net17 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP2 Z B net016 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 net016 net17 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 AN VDD VSS net17 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR2BX0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2BX0P7H7L AN B VDD VSS Z
*.PININFO AN:I B:I Z:O VDD:B VSS:B
MMN2 Z B VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN0 Z net17 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMP2 Z B net016 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP1 net016 net17 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
XXI3 AN VDD VSS net17 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR2BX12H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2BX12H7L AN B VDD VSS Z
*.PININFO AN:I B:I Z:O VDD:B VSS:B
MMN2 Z B VSS VSS nm1p2_lvt_lp W=1.8u L=60n m=1
MMN0 Z net17 VSS VSS nm1p2_lvt_lp W=1.8u L=60n m=1
MMP2 Z B net016 VDD pm1p2_lvt_lp W=2.28u L=60n m=1
MMP1 net016 net17 VDD VDD pm1p2_lvt_lp W=2.28u L=60n m=1
XXI3 AN VDD VSS net17 / INV pl=6e-08 pw=7.6e-07 nl=6e-08 nw=6e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR2BX16H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2BX16H7L AN B VDD VSS Z
*.PININFO AN:I B:I Z:O VDD:B VSS:B
MMN2 Z B VSS VSS nm1p2_lvt_lp W=2.4u L=60n m=1
MMN0 Z net17 VSS VSS nm1p2_lvt_lp W=2.4u L=60n m=1
MMP2 Z B net016 VDD pm1p2_lvt_lp W=3.04u L=60n m=1
MMP1 net016 net17 VDD VDD pm1p2_lvt_lp W=3.04u L=60n m=1
XXI3 AN VDD VSS net17 / INV pl=6e-08 pw=11.4e-07 nl=6e-08 nw=9e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR2BX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2BX1H7L AN B VDD VSS Z
*.PININFO AN:I B:I Z:O VDD:B VSS:B
MMN2 Z B VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN0 Z net17 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMP2 Z B net016 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP1 net016 net17 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
XXI3 AN VDD VSS net17 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR2BX1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2BX1P4H7L AN B VDD VSS Z
*.PININFO AN:I B:I Z:O VDD:B VSS:B
MMN2 Z B VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN0 Z net17 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMP2 Z B net016 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP1 net016 net17 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
XXI3 AN VDD VSS net17 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR2BX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2BX2H7L AN B VDD VSS Z
*.PININFO AN:I B:I Z:O VDD:B VSS:B
MMN2 Z B VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN0 Z net17 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP2 Z B net016 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP1 net016 net17 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
XXI3 AN VDD VSS net17 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR2BX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2BX3H7L AN B VDD VSS Z
*.PININFO AN:I B:I Z:O VDD:B VSS:B
MMN2 Z B VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN0 Z net17 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMP2 Z B net016 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP1 net016 net17 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
XXI3 AN VDD VSS net17 / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR2BX4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2BX4H7L AN B VDD VSS Z
*.PININFO AN:I B:I Z:O VDD:B VSS:B
MMN2 Z B VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN0 Z net17 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMP2 Z B net016 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP1 net016 net17 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
XXI3 AN VDD VSS net17 / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR2BX6H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2BX6H7L AN B VDD VSS Z
*.PININFO AN:I B:I Z:O VDD:B VSS:B
MMN2 Z B VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN0 Z net17 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMP2 Z B net016 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP1 net016 net17 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
XXI3 AN VDD VSS net17 / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR2BX8H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2BX8H7L AN B VDD VSS Z
*.PININFO AN:I B:I Z:O VDD:B VSS:B
MMN2 Z B VSS VSS nm1p2_lvt_lp W=1.2u L=60n m=1
MMN0 Z net17 VSS VSS nm1p2_lvt_lp W=1.2u L=60n m=1
MMP2 Z B net016 VDD pm1p2_lvt_lp W=1.52u L=60n m=1
MMP1 net016 net17 VDD VDD pm1p2_lvt_lp W=1.52u L=60n m=1
XXI3 AN VDD VSS net17 / INV pl=6e-08 pw=6.2e-07 nl=6e-08 nw=5e-07
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR2X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2X0P5H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MNM0 Y B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 Y A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM0 Y B net015 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 net015 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR2X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2X0P7H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MNM0 Y B VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN0 Y A VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MPM0 Y B net015 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP1 net015 A VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR2X12H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2X12H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MNM0 Y B VSS VSS nm1p2_lvt_lp W=1.8u L=60n m=1
MMN0 Y A VSS VSS nm1p2_lvt_lp W=1.8u L=60n m=1
MPM0 Y B net015 VDD pm1p2_lvt_lp W=2.28u L=60n m=1
MMP1 net015 A VDD VDD pm1p2_lvt_lp W=2.28u L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR2X16H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2X16H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MNM0 Y B VSS VSS nm1p2_lvt_lp W=2.4u L=60n m=1
MMN0 Y A VSS VSS nm1p2_lvt_lp W=2.4u L=60n m=1
MPM0 Y B net015 VDD pm1p2_lvt_lp W=3.04u L=60n m=1
MMP1 net015 A VDD VDD pm1p2_lvt_lp W=3.04u L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR2X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2X1H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MNM0 Y B VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN0 Y A VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MPM0 Y B net015 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP1 net015 A VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR2X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2X1P4H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MNM0 Y B VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN0 Y A VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MPM0 Y B net015 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP1 net015 A VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR2X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2X2H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MNM0 Y B VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN0 Y A VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MPM0 Y B net015 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP1 net015 A VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR2X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2X3H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MNM0 Y B VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN0 Y A VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MPM0 Y B net015 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP1 net015 A VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR2X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2X4H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MNM0 Y B VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN0 Y A VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MPM0 Y B net015 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP1 net015 A VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR2X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2X6H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MNM0 Y B VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN0 Y A VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MPM0 Y B net015 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP1 net015 A VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR2X8H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2X8H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MNM0 Y B VSS VSS nm1p2_lvt_lp W=1.2u L=60n m=1
MMN0 Y A VSS VSS nm1p2_lvt_lp W=1.2u L=60n m=1
MPM0 Y B net015 VDD pm1p2_lvt_lp W=1.52u L=60n m=1
MMP1 net015 A VDD VDD pm1p2_lvt_lp W=1.52u L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR3BX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR3BX0P5H7L AN B C VDD VSS Y
*.PININFO AN:I B:I C:I Y:O VDD:B VSS:B
MMN3 Y net17 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 Y C VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 Y B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP3 Y C net026 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 net020 net17 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP2 net026 B net020 VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 AN VDD VSS net17 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR3BX0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR3BX0P7H7L AN B C VDD VSS Y
*.PININFO AN:I B:I C:I Y:O VDD:B VSS:B
MMN3 Y net17 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN2 Y C VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN0 Y B VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMP3 Y C net026 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP1 net020 net17 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP2 net026 B net020 VDD pm1p2_lvt_lp W=222n L=60n m=1
XXI3 AN VDD VSS net17 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR3BX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR3BX1H7L AN B C VDD VSS Y
*.PININFO AN:I B:I C:I Y:O VDD:B VSS:B
MMN3 Y net17 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN2 Y C VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN0 Y B VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMP3 Y C net026 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP1 net020 net17 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP2 net026 B net020 VDD pm1p2_lvt_lp W=270n L=60n m=1
XXI3 AN VDD VSS net17 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR3BX1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR3BX1P4H7L AN B C VDD VSS Y
*.PININFO AN:I B:I C:I Y:O VDD:B VSS:B
MMN3 Y net17 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN2 Y C VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN0 Y B VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMP3 Y C net026 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP1 net020 net17 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP2 net026 B net020 VDD pm1p2_lvt_lp W=314n L=60n m=1
XXI3 AN VDD VSS net17 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR3BX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR3BX2H7L AN B C VDD VSS Y
*.PININFO AN:I B:I C:I Y:O VDD:B VSS:B
MMN3 Y net17 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN2 Y C VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN0 Y B VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP3 Y C net026 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP1 net020 net17 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP2 net026 B net020 VDD pm1p2_lvt_lp W=380n L=60n m=1
XXI3 AN VDD VSS net17 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR3BX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR3BX3H7L AN B C VDD VSS Y
*.PININFO AN:I B:I C:I Y:O VDD:B VSS:B
MMN3 Y net17 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN2 Y C VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN0 Y B VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMP3 Y C net026 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP1 net020 net17 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP2 net026 B net020 VDD pm1p2_lvt_lp W=570n L=60n m=1
XXI3 AN VDD VSS net17 / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR3BX4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR3BX4H7L AN B C VDD VSS Y
*.PININFO AN:I B:I C:I Y:O VDD:B VSS:B
MMN3 Y net17 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN2 Y C VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN0 Y B VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMP3 Y C net026 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP1 net020 net17 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP2 net026 B net020 VDD pm1p2_lvt_lp W=760n L=60n m=1
XXI3 AN VDD VSS net17 / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR3BX6H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR3BX6H7L AN B C VDD VSS Y
*.PININFO AN:I B:I C:I Y:O VDD:B VSS:B
MMN3 Y net17 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN2 Y C VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN0 Y B VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMP3 Y C net026 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP1 net020 net17 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP2 net026 B net020 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
XXI3 AN VDD VSS net17 / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR3X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR3X0P5H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN3 Y A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 Y C VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 Y B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP3 Y C net025 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 net019 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP2 net025 B net019 VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR3X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR3X0P7H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN3 Y A VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN2 Y C VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN0 Y B VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMP3 Y C net025 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP1 net019 A VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP2 net025 B net019 VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR3X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR3X1H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN3 Y A VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN2 Y C VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN0 Y B VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMP3 Y C net025 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP1 net019 A VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP2 net025 B net019 VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR3X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR3X1P4H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN3 Y A VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN2 Y C VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN0 Y B VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMP3 Y C net025 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP1 net019 A VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP2 net025 B net019 VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR3X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR3X2H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN3 Y A VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN2 Y C VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN0 Y B VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP3 Y C net025 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP1 net019 A VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP2 net025 B net019 VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR3X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR3X3H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN3 Y A VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN2 Y C VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN0 Y B VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMP3 Y C net025 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP1 net019 A VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP2 net025 B net019 VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR3X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR3X4H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN3 Y A VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN2 Y C VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN0 Y B VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMP3 Y C net025 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP1 net019 A VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP2 net025 B net019 VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR3X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR3X6H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN3 Y A VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN2 Y C VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN0 Y B VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMP3 Y C net025 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP1 net019 A VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP2 net025 B net019 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR3X8H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR3X8H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MMN3 Y A VSS VSS nm1p2_lvt_lp W=1.2u L=60n m=1
MMN2 Y C VSS VSS nm1p2_lvt_lp W=1.2u L=60n m=1
MMN0 Y B VSS VSS nm1p2_lvt_lp W=1.2u L=60n m=1
MMP3 Y C net025 VDD pm1p2_lvt_lp W=1.52u L=60n m=1
MMP1 net019 A VDD VDD pm1p2_lvt_lp W=1.52u L=60n m=1
MMP2 net025 B net019 VDD pm1p2_lvt_lp W=1.52u L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR4BBX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4BBX0P5H7L AN BN C D VDD VSS Y
*.PININFO AN:I BN:I C:I D:I Y:O VDD:B VSS:B
MMN4 Y net17 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN3 Y net47 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 Y D VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 Y C VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP4 Y D net27 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP3 net27 C net031 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 net025 net17 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP2 net031 net47 net025 VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI0 BN VDD VSS net47 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XI1 AN VDD VSS net17 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR4BBX0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4BBX0P7H7L AN BN C D VDD VSS Y
*.PININFO AN:I BN:I C:I D:I Y:O VDD:B VSS:B
MMN4 Y net17 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN3 Y net47 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN2 Y D VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN0 Y C VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMP4 Y D net27 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP3 net27 C net031 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP1 net025 net17 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP2 net031 net47 net025 VDD pm1p2_lvt_lp W=222n L=60n m=1
XI1 AN VDD VSS net17 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI0 BN VDD VSS net47 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR4BBX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4BBX1H7L AN BN C D VDD VSS Y
*.PININFO AN:I BN:I C:I D:I Y:O VDD:B VSS:B
MMN4 Y net17 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN3 Y net47 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN2 Y D VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN0 Y C VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMP4 Y D net27 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP3 net27 C net031 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP1 net025 net17 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP2 net031 net47 net025 VDD pm1p2_lvt_lp W=270n L=60n m=1
XI1 AN VDD VSS net17 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI0 BN VDD VSS net47 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR4BBX1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4BBX1P4H7L AN BN C D VDD VSS Y
*.PININFO AN:I BN:I C:I D:I Y:O VDD:B VSS:B
MMN4 Y net17 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN3 Y net47 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN2 Y D VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN0 Y C VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMP4 Y D net27 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP3 net27 C net031 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP1 net025 net17 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP2 net031 net47 net025 VDD pm1p2_lvt_lp W=314n L=60n m=1
XI1 AN VDD VSS net17 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI0 BN VDD VSS net47 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR4BBX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4BBX2H7L AN BN C D VDD VSS Y
*.PININFO AN:I BN:I C:I D:I Y:O VDD:B VSS:B
MMN4 Y net17 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN3 Y net47 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN2 Y D VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN0 Y C VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP4 Y D net27 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP3 net27 C net031 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP1 net025 net17 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP2 net031 net47 net025 VDD pm1p2_lvt_lp W=380n L=60n m=1
XI1 AN VDD VSS net17 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI0 BN VDD VSS net47 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR4BBX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4BBX3H7L AN BN C D VDD VSS Y
*.PININFO AN:I BN:I C:I D:I Y:O VDD:B VSS:B
MMN4 Y net17 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN3 Y net47 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN2 Y D VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN0 Y C VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMP4 Y D net27 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP3 net27 C net031 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP1 net025 net17 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP2 net031 net47 net025 VDD pm1p2_lvt_lp W=570n L=60n m=1
XXI5 BN VDD VSS net47 / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
XI2 AN VDD VSS net17 / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR4BBX4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4BBX4H7L AN BN C D VDD VSS Y
*.PININFO AN:I BN:I C:I D:I Y:O VDD:B VSS:B
MMN4 Y net17 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN3 Y net47 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN2 Y D VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN0 Y C VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMP4 Y D net27 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP3 net27 C net031 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP1 net025 net17 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP2 net031 net47 net025 VDD pm1p2_lvt_lp W=760n L=60n m=1
XI3 BN VDD VSS net47 / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
XI2 AN VDD VSS net17 / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR4BX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4BX0P5H7L AN B C D VDD VSS Y
*.PININFO AN:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 Y net17 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN3 Y B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 Y D VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 Y C VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP4 Y D net27 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP3 net27 C net030 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 net024 net17 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP2 net030 B net024 VDD pm1p2_lvt_lp W=190n L=60n m=1
XI1 AN VDD VSS net17 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR4BX0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4BX0P7H7L AN B C D VDD VSS Y
*.PININFO AN:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 Y net17 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN3 Y B VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN2 Y D VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN0 Y C VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMP4 Y D net27 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP3 net27 C net030 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP1 net024 net17 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP2 net030 B net024 VDD pm1p2_lvt_lp W=222n L=60n m=1
XI1 AN VDD VSS net17 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR4BX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4BX1H7L AN B C D VDD VSS Y
*.PININFO AN:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 Y net17 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN3 Y B VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN2 Y D VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN0 Y C VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMP4 Y D net27 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP3 net27 C net030 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP1 net024 net17 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP2 net030 B net024 VDD pm1p2_lvt_lp W=270n L=60n m=1
XI1 AN VDD VSS net17 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR4BX1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4BX1P4H7L AN B C D VDD VSS Z
*.PININFO AN:I B:I C:I D:I Z:O VDD:B VSS:B
MMN4 Z net17 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN3 Z B VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN2 Z D VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN0 Z C VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMP4 Z D net27 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP3 net27 C net030 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP1 net024 net17 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP2 net030 B net024 VDD pm1p2_lvt_lp W=314n L=60n m=1
XI1 AN VDD VSS net17 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR4BX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4BX2H7L AN B C D VDD VSS Y
*.PININFO AN:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 Y net17 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN3 Y B VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN2 Y D VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN0 Y C VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP4 Y D net27 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP3 net27 C net030 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP1 net024 net17 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP2 net030 B net024 VDD pm1p2_lvt_lp W=380n L=60n m=1
XI1 AN VDD VSS net17 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR4BX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4BX3H7L AN B C D VDD VSS Y
*.PININFO AN:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 Y net17 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN3 Y B VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN2 Y D VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN0 Y C VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMP4 Y D net27 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP3 net27 C net030 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP1 net024 net17 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP2 net030 B net024 VDD pm1p2_lvt_lp W=570n L=60n m=1
XXI3 AN VDD VSS net17 / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR4BX4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4BX4H7L AN B C D VDD VSS Y
*.PININFO AN:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 Y net17 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN3 Y B VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN2 Y D VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN0 Y C VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMP4 Y D net27 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP3 net27 C net030 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP1 net024 net17 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP2 net030 B net024 VDD pm1p2_lvt_lp W=760n L=60n m=1
XXI3 AN VDD VSS net17 / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR4X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4X0P5H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 Y A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN3 Y B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 Y D VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 Y C VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP4 Y D net27 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP3 net27 C net029 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 net023 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP2 net029 B net023 VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR4X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4X0P7H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 Y A VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN3 Y B VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN2 Y D VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN0 Y C VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMP4 Y D net27 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP3 net27 C net029 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP1 net023 A VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP2 net029 B net023 VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR4X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4X1H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 Y A VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN3 Y B VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN2 Y D VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN0 Y C VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMP4 Y D net27 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP3 net27 C net029 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP1 net023 A VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP2 net029 B net023 VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR4X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4X1P4H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 Y A VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN3 Y B VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN2 Y D VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN0 Y C VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMP4 Y D net27 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP3 net27 C net029 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP1 net023 A VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP2 net029 B net023 VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR4X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4X2H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 Y A VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN3 Y B VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN2 Y D VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN0 Y C VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP4 Y D net27 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP3 net27 C net029 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP1 net023 A VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP2 net029 B net023 VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR4X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4X3H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 Y A VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN3 Y B VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN2 Y D VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN0 Y C VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMP4 Y D net27 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP3 net27 C net029 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP1 net023 A VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP2 net029 B net023 VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR4X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4X4H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 Y A VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN3 Y B VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN2 Y D VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN0 Y C VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMP4 Y D net27 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP3 net27 C net029 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP1 net023 A VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP2 net029 B net023 VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    NOR4X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4X6H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MMN4 Y A VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN3 Y B VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN2 Y D VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN0 Y C VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMP4 Y D net27 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP3 net27 C net029 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP1 net023 A VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP2 net029 B net023 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA211X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA211X0P5H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 net10 C0 net30 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 net22 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net22 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net30 B0 net22 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM1 net10 A1 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 net10 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM2 net10 C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net10 VDD VSS Y / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA211X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA211X0P7H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 net10 C0 net30 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 net22 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net22 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net30 B0 net22 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM1 net10 A1 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 net10 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM2 net10 C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net10 VDD VSS Y / INV pl=6e-08 pw=2.22e-07 nl=6e-08 nw=1.74e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA211X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA211X1H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 net10 C0 net30 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 net22 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net22 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net30 B0 net22 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM1 net10 A1 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 net10 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM2 net10 C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net10 VDD VSS Y / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA211X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA211X1P4H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 net10 C0 net30 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 net22 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net22 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net30 B0 net22 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM1 net10 A1 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 net10 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM2 net10 C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net10 VDD VSS Y / INV pl=6e-08 pw=3.14e-07 nl=6e-08 nw=2.46e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA211X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA211X2H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 net10 C0 net30 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 net22 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net22 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net30 B0 net22 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM1 net10 A1 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 net10 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM2 net10 C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net10 VDD VSS Y / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA211X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA211X3H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 net10 C0 net30 VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM4 net22 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM3 net30 B0 net22 VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM5 net22 A1 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMPM1 net10 A1 net13 VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM5 net10 C0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM3 net13 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM4 net10 B0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
XXI3 net10 VDD VSS Y / INV pl=6e-08 pw=5.7e-07 nl=6e-08 nw=4.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA211X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA211X4H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 net10 C0 net30 VSS nm1p2_lvt_lp W=250n L=60n m=1
MNM4 net22 A0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MNM3 net30 B0 net22 VSS nm1p2_lvt_lp W=250n L=60n m=1
MNM5 net22 A1 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMPM1 net10 A1 net13 VDD pm1p2_lvt_lp W=310n L=60n m=1
MPM5 net10 C0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MPM3 net13 A0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MPM4 net10 B0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
XXI3 net10 VDD VSS Y / INV pl=6e-08 pw=7.6e-07 nl=6e-08 nw=6e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA211X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA211X6H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 net10 C0 net30 VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM4 net22 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM3 net30 B0 net22 VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM5 net22 A1 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMPM1 net10 A1 net13 VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM5 net10 C0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM3 net13 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM4 net10 B0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
XXI3 net10 VDD VSS Y / INV pl=6e-08 pw=11.4e-07 nl=6e-08 nw=9e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA21X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA21X0P5H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMNM2 net11 B0 net27 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net27 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net27 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM1 net11 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net11 A1 net14 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net14 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net11 VDD VSS Y / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA21X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA21X0P7H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMNM2 net11 B0 net27 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net27 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net27 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM1 net11 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net11 A1 net14 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net14 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net11 VDD VSS Y / INV pl=6e-08 pw=2.22e-07 nl=6e-08 nw=1.74e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA21X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA21X1H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MNM0 net27 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net27 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net_04 B0 net27 VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM0 net_04 A1 net14 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM2 net14 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM3 net_04 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net_04 VDD VSS Y / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA21X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA21X1P4H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMNM2 net11 B0 net27 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net27 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net27 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM1 net11 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net11 A1 net14 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net14 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net11 VDD VSS Y / INV pl=6e-08 pw=3.14e-07 nl=6e-08 nw=2.46e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA21X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA21X2H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMNM2 net11 B0 net27 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net27 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net27 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM1 net11 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net11 A1 net14 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net14 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net11 VDD VSS Y / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA21X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA21X3H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMNM2 net11 B0 net27 VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM0 net27 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM1 net27 A1 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MPM1 net11 B0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM0 net11 A1 net14 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM0 net14 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
XXI3 net11 VDD VSS Y / INV pl=6e-08 pw=5.7e-07 nl=6e-08 nw=4.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA21X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA21X4H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMNM2 net11 B0 net27 VSS nm1p2_lvt_lp W=250n L=60n m=1
MNM0 net27 A0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MNM1 net27 A1 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MPM1 net11 B0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MPM0 net11 A1 net14 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM0 net14 A0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
XXI3 net11 VDD VSS Y / INV pl=6e-08 pw=7.6e-07 nl=6e-08 nw=6e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA21X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA21X6H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMNM2 net11 B0 net27 VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM0 net27 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM1 net27 A1 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MPM1 net11 B0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM0 net11 A1 net14 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM0 net14 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
XXI3 net11 VDD VSS Y / INV pl=6e-08 pw=11.4e-07 nl=6e-08 nw=9e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA21X8H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA21X8H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MMNM2 net11 B0 net27 VSS nm1p2_lvt_lp W=500n L=60n m=1
MNM0 net27 A0 VSS VSS nm1p2_lvt_lp W=500n L=60n m=1
MNM1 net27 A1 VSS VSS nm1p2_lvt_lp W=500n L=60n m=1
MPM1 net11 B0 VDD VDD pm1p2_lvt_lp W=620n L=60n m=1
MPM0 net11 A1 net14 VDD pm1p2_lvt_lp W=620n L=60n m=1
MMPM0 net14 A0 VDD VDD pm1p2_lvt_lp W=620n L=60n m=1
XXI3 net11 VDD VSS Y / INV pl=6e-08 pw=15.2e-07 nl=6e-08 nw=12e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA221X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA221X0P5H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MNM3 net15 C0 net31 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net31 B0 net39 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 net31 B1 net39 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net39 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net39 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM1 net22 B1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net18 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM3 net15 C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net15 A0 net18 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM2 net15 B0 net22 VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net15 VDD VSS Y / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA221X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA221X0P7H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MNM3 net15 C0 net31 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net31 B0 net39 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 net31 B1 net39 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net39 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net39 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM1 net22 B1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net18 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM3 net15 C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net15 A0 net18 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM2 net15 B0 net22 VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net15 VDD VSS Y / INV pl=6e-08 pw=2.22e-07 nl=6e-08 nw=1.74e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA221X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA221X1H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MNM6 net31 B0 net39 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM5 net31 B1 net39 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM4 net39 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM7 net15 C0 net31 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net39 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM4 net15 B0 net22 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net15 A0 net18 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM7 net15 C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM6 net18 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM5 net22 B1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net15 VDD VSS Y / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA221X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA221X1P4H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MNM3 net15 C0 net31 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net31 B0 net39 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 net31 B1 net39 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net39 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net39 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM1 net22 B1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net18 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM3 net15 C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net15 A0 net18 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM2 net15 B0 net22 VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net15 VDD VSS Y / INV pl=6e-08 pw=3.14e-07 nl=6e-08 nw=2.46e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA221X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA221X2H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MNM3 net15 C0 net31 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net31 B0 net39 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 net31 B1 net39 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net39 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net39 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM1 net22 B1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net18 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM3 net15 C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net15 A0 net18 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM2 net15 B0 net22 VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net15 VDD VSS Y / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA221X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA221X3H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MNM3 net15 C0 net31 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM3 net31 B0 net39 VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM2 net31 B1 net39 VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM0 net39 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM1 net39 A1 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MPM1 net22 B1 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM0 net18 A1 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM3 net15 C0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM1 net15 A0 net18 VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM2 net15 B0 net22 VDD pm1p2_lvt_lp W=270n L=60n m=1
XXI1 net15 VDD VSS Y / INV pl=6e-08 pw=5.7e-07 nl=6e-08 nw=4.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA221X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA221X4H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MNM3 net15 C0 net31 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM3 net31 B0 net39 VSS nm1p2_lvt_lp W=250n L=60n m=1
MNM2 net31 B1 net39 VSS nm1p2_lvt_lp W=250n L=60n m=1
MNM0 net39 A0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MNM1 net39 A1 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MPM1 net22 B1 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MPM0 net18 A1 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MPM3 net15 C0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM1 net15 A0 net18 VDD pm1p2_lvt_lp W=310n L=60n m=1
MPM2 net15 B0 net22 VDD pm1p2_lvt_lp W=310n L=60n m=1
XXI1 net15 VDD VSS Y / INV pl=6e-08 pw=7.6e-07 nl=6e-08 nw=6e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA222X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA222X0P5H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 net082 C1 net44 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM4 net082 C0 net44 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net44 B1 net52 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net44 B0 net52 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net52 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net52 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM5 net082 C1 net11 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM4 net11 C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net082 B1 net19 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net19 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net082 A1 net27 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net27 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net082 VDD VSS Y / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA222X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA222X0P7H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 net082 C1 net44 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM4 net082 C0 net44 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net44 B1 net52 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net44 B0 net52 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net52 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net52 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM5 net082 C1 net11 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM4 net11 C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net082 B1 net19 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net19 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net082 A1 net27 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net27 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net082 VDD VSS Y / INV pl=6e-08 pw=2.22e-07 nl=6e-08 nw=1.74e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA222X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA222X1H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 net082 C1 net44 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM4 net082 C0 net44 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net44 B1 net52 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net44 B0 net52 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net52 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net52 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM5 net082 C1 net11 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM4 net11 C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net082 B1 net19 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net19 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net082 A1 net27 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net27 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net082 VDD VSS Y / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA222X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA222X1P4H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 net082 C1 net44 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM4 net082 C0 net44 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net44 B1 net52 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net44 B0 net52 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net52 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net52 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM5 net082 C1 net11 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM4 net11 C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net082 B1 net19 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net19 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net082 A1 net27 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net27 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net082 VDD VSS Y / INV pl=6e-08 pw=3.14e-07 nl=6e-08 nw=2.46e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA222X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA222X2H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 net082 C1 net44 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM4 net082 C0 net44 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net44 B1 net52 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net44 B0 net52 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net52 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net52 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM5 net082 C1 net11 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM4 net11 C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net082 B1 net19 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net19 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net082 A1 net27 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net27 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net082 VDD VSS Y / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA222X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA222X3H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 net082 C1 net44 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM4 net082 C0 net44 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM3 net44 B1 net52 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM2 net44 B0 net52 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM1 net52 A1 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM0 net52 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMPM5 net082 C1 net11 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM4 net11 C0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM3 net082 B1 net19 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM2 net19 B0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM1 net082 A1 net27 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM0 net27 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
XXI3 net082 VDD VSS Y / INV pl=6e-08 pw=5.7e-07 nl=6e-08 nw=4.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA222X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA222X4H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 net082 C1 net44 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM4 net082 C0 net44 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM3 net44 B1 net52 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM2 net44 B0 net52 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM1 net52 A1 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM0 net52 A0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMPM5 net082 C1 net11 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM4 net11 C0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM3 net082 B1 net19 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM2 net19 B0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM1 net082 A1 net27 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM0 net27 A0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
XXI3 net082 VDD VSS Y / INV pl=6e-08 pw=7.6e-07 nl=6e-08 nw=6e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA22X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA22X0P5H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MNM2 net34 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net10 B0 net34 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net34 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net10 B1 net34 VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM1 net10 B1 net21 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net10 A1 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net13 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM2 net21 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net10 VDD VSS Y / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA22X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA22X0P7H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MNM2 net34 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net10 B0 net34 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net34 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net10 B1 net34 VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM1 net10 B1 net21 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net10 A1 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net13 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM2 net21 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net10 VDD VSS Y / INV pl=6e-08 pw=2.22e-07 nl=6e-08 nw=1.74e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA22X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA22X1H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MNM1 net34 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 net34 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM3 net10 B1 net34 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net10 B0 net34 VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM3 net10 B1 net21 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM2 net21 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 S A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net10 A1 S VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net10 VDD VSS Y / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA22X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA22X1P4H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MNM2 net34 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net10 B0 net34 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net34 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net10 B1 net34 VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM1 net10 B1 net21 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net10 A1 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net13 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM2 net21 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net10 VDD VSS Y / INV pl=6e-08 pw=3.14e-07 nl=6e-08 nw=2.46e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA22X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA22X2H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MNM0 net10 B0 net34 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 net34 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM3 net34 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net10 B1 net34 VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM3 net21 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM2 net13 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 net10 B1 net21 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net10 A1 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI1 net10 VDD VSS Y / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA22X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA22X3H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MNM0 net10 B0 net34 VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM3 net34 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM2 net34 A1 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM1 net10 B1 net34 VSS nm1p2_lvt_lp W=210n L=60n m=1
MPM1 net10 B1 net21 VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM2 net13 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM3 net21 B0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM0 net10 A1 net13 VDD pm1p2_lvt_lp W=270n L=60n m=1
XXI1 net10 VDD VSS Y / INV pl=6e-08 pw=5.7e-07 nl=6e-08 nw=4.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA22X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA22X4H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MNM0 net10 B0 net34 VSS nm1p2_lvt_lp W=250n L=60n m=1
MNM3 net34 A0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MNM2 net34 A1 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MNM1 net10 B1 net34 VSS nm1p2_lvt_lp W=250n L=60n m=1
MPM1 net10 B1 net21 VDD pm1p2_lvt_lp W=310n L=60n m=1
MPM2 net13 A0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MPM3 net21 B0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MPM0 net10 A1 net13 VDD pm1p2_lvt_lp W=310n L=60n m=1
XXI1 net10 VDD VSS Y / INV pl=6e-08 pw=7.6e-07 nl=6e-08 nw=6e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA22X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA22X6H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MNM0 net10 B0 net34 VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM3 net34 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM2 net34 A1 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM1 net10 B1 net34 VSS nm1p2_lvt_lp W=300n L=60n m=1
MPM1 net10 B1 net21 VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM2 net13 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM3 net21 B0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM0 net10 A1 net13 VDD pm1p2_lvt_lp W=380n L=60n m=1
XXI1 net10 VDD VSS Y / INV pl=6e-08 pw=11.4e-07 nl=6e-08 nw=9e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA31X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA31X0P5H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMNM3 net045 B0 net34 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net34 A2 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net34 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net34 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM2 net17 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net045 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 net13 A1 net17 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net045 A2 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net045 VDD VSS Y / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA31X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA31X0P7H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMNM3 net045 B0 net34 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net34 A2 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net34 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net34 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM2 net17 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net045 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 net13 A1 net17 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net045 A2 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net045 VDD VSS Y / INV pl=6e-08 pw=2.22e-07 nl=6e-08 nw=1.74e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA31X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA31X1H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMNM3 net045 B0 net34 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net34 A2 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net34 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net34 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM2 net17 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net045 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 net13 A1 net17 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net045 A2 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net045 VDD VSS Y / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA31X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA31X1P4H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMNM3 net045 B0 net34 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net34 A2 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net34 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net34 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM2 net17 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net045 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 net13 A1 net17 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net045 A2 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net045 VDD VSS Y / INV pl=6e-08 pw=3.14e-07 nl=6e-08 nw=2.46e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA31X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA31X2H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMNM3 net045 B0 net34 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net34 A2 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net34 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net34 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM2 net17 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net045 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 net13 A1 net17 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net045 A2 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 net045 VDD VSS Y / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA31X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA31X3H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMNM3 net045 B0 net34 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM2 net34 A2 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM1 net34 A1 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM0 net34 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MPM2 net17 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM3 net045 B0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM1 net13 A1 net17 VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM0 net045 A2 net13 VDD pm1p2_lvt_lp W=270n L=60n m=1
XXI3 net045 VDD VSS Y / INV pl=6e-08 pw=5.7e-07 nl=6e-08 nw=4.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OA31X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OA31X4H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMNM3 net045 B0 net34 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM2 net34 A2 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM1 net34 A1 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM0 net34 A0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MPM2 net17 A0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM3 net045 B0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MPM1 net13 A1 net17 VDD pm1p2_lvt_lp W=310n L=60n m=1
MPM0 net045 A2 net13 VDD pm1p2_lvt_lp W=310n L=60n m=1
XXI3 net045 VDD VSS Y / INV pl=6e-08 pw=7.6e-07 nl=6e-08 nw=6e-07
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI211X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI211X0P5H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 Y C0 net30 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 net22 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net22 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net30 B0 net22 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM1 Y A1 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 Y B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM2 Y C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI211X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI211X0P7H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 Y C0 net30 VSS nm1p2_lvt_lp W=175n L=60n m=1
MNM2 net22 A1 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MNM1 net22 A0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MNM0 net30 B0 net22 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMPM1 Y A1 net13 VDD pm1p2_lvt_lp W=222n L=60n m=1
MPM1 Y B0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MPM2 Y C0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI211X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI211X1H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 Y C0 net30 VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM4 net22 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM3 net30 B0 net22 VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM5 net22 A1 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MPM5 Y C0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM4 Y B0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM3 Y A1 net13 VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI211X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI211X1P4H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 Y C0 net30 VSS nm1p2_lvt_lp W=245n L=60n m=1
MNM2 net22 A1 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MNM1 net22 A0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MNM0 net30 B0 net22 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMPM1 Y A1 net13 VDD pm1p2_lvt_lp W=314n L=60n m=1
MPM1 Y B0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MPM2 Y C0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI211X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI211X2H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 Y C0 net30 VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM4 net22 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM3 net30 B0 net22 VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM5 net22 A1 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMPM1 Y A1 net13 VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM5 Y C0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM3 net13 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM4 Y B0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI211X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI211X3H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 Y C0 net30 VSS nm1p2_lvt_lp W=450n L=60n m=1
MNM2 net22 A1 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MNM1 net22 A0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MNM0 net30 B0 net22 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMPM1 Y A1 net13 VDD pm1p2_lvt_lp W=570n L=60n m=1
MPM1 Y B0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MPM2 Y C0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI211X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI211X4H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MNM7 net22 A0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MNM8 net22 A1 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MNM6 net30 B0 net22 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM3 Y C0 net30 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMPM1 Y A1 net13 VDD pm1p2_lvt_lp W=760n L=60n m=1
MPM7 Y C0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MPM8 net13 A0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MPM6 Y B0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI211X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI211X6H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMNM3 Y C0 net30 VSS nm1p2_lvt_lp W=900n L=60n m=1
MNM2 net22 A1 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MNM1 net22 A0 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MNM0 net30 B0 net22 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMPM1 Y A1 net13 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MPM1 Y B0 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MPM2 Y C0 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI21BX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI21BX0P5H7L A0 A1 B0N VDD VSS Y
*.PININFO A0:I A1:I B0N:I Y:O VDD:B VSS:B
MMNM2 Y net30 net17 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net17 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net17 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM1 Y A1 net12 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 Y net30 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net12 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI0 B0N VDD VSS net30 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI21BX0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI21BX0P7H7L A0 A1 B0N VDD VSS Y
*.PININFO A0:I A1:I B0N:I Y:O VDD:B VSS:B
MMNM2 Y net30 net17 VSS nm1p2_lvt_lp W=175n L=60n m=1
MNM0 net17 A0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MNM1 net17 A1 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MPM1 Y A1 net12 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM2 Y net30 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MPM0 net12 A0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
XXI0 B0N VDD VSS net30 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI21BX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI21BX1H7L A0 A1 B0N VDD VSS Y
*.PININFO A0:I A1:I B0N:I Y:O VDD:B VSS:B
MNM0 net17 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM1 net17 A1 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM2 Y net30 net17 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMPM2 Y net30 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM0 Y A1 net12 VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM1 net12 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
XXI0 B0N VDD VSS net30 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI21BX1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI21BX1P4H7L A0 A1 B0N VDD VSS Y
*.PININFO A0:I A1:I B0N:I Y:O VDD:B VSS:B
MMNM2 Y net30 net17 VSS nm1p2_lvt_lp W=245n L=60n m=1
MNM0 net17 A0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MNM1 net17 A1 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MPM1 Y A1 net12 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM2 Y net30 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MPM0 net12 A0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
XXI0 B0N VDD VSS net30 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI21BX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI21BX2H7L A0 A1 B0N VDD VSS Y
*.PININFO A0:I A1:I B0N:I Y:O VDD:B VSS:B
MMNM2 Y net30 net17 VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM1 net17 A1 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM0 net17 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MPM1 Y A1 net12 VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM2 net12 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM0 Y net30 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
XXI0 B0N VDD VSS net30 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI21BX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI21BX3H7L A0 A1 B0N VDD VSS Y
*.PININFO A0:I A1:I B0N:I Y:O VDD:B VSS:B
MNM0 Y net30 net17 VSS nm1p2_lvt_lp W=450n L=60n m=1
MNM2 net17 A1 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MNM1 net17 A0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MPM1 Y A1 net12 VDD pm1p2_lvt_lp W=570n L=60n m=1
MPM2 net12 A0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MPM0 Y net30 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
XXI0 B0N VDD VSS net30 / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI21BX4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI21BX4H7L A0 A1 B0N VDD VSS Y
*.PININFO A0:I A1:I B0N:I Y:O VDD:B VSS:B
MNM0 Y net30 net17 VSS nm1p2_lvt_lp W=600n L=60n m=1
MNM2 net17 A1 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MNM1 net17 A0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MPM1 Y A1 net12 VDD pm1p2_lvt_lp W=760n L=60n m=1
MPM2 net12 A0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MPM0 Y net30 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
XXI0 B0N VDD VSS net30 / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI21BX6H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI21BX6H7L A0 A1 B0N VDD VSS Y
*.PININFO A0:I A1:I B0N:I Y:O VDD:B VSS:B
MNM0 Y net30 net17 VSS nm1p2_lvt_lp W=900n L=60n m=1
MNM2 net17 A1 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MNM1 net17 A0 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MPM1 Y A1 net12 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MPM2 net12 A0 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MPM0 Y net30 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
XXI0 B0N VDD VSS net30 / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI21X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI21X0P5H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MNM1 net8 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 Y B0 net8 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net8 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM1 Y B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP3 net033 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 Y A1 net033 VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI21X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI21X0P7H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MNM1 net8 A1 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN5 Y B0 net8 VSS nm1p2_lvt_lp W=175n L=60n m=1
MNM0 net8 A0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MPM1 Y B0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP3 net033 A0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MPM0 Y A1 net033 VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI21X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI21X1H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MNM1 net8 A1 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN5 Y B0 net8 VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM0 net8 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MPM0 Y A1 net033 VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM1 net033 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP4 Y B0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI21X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI21X1P4H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MNM1 net8 A1 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN5 Y B0 net8 VSS nm1p2_lvt_lp W=245n L=60n m=1
MNM0 net8 A0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MPM1 Y B0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP3 net033 A0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MPM0 Y A1 net033 VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI21X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI21X2H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MNM1 net8 A1 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM0 net8 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN5 Y B0 net8 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP3 net033 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM1 Y B0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM0 Y A1 net033 VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI21X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI21X3H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MNM1 net8 A1 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MNM0 net8 A0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN5 Y B0 net8 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMP3 net033 A0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MPM1 Y B0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MPM0 Y A1 net033 VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI21X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI21X4H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MNM1 net8 A1 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MNM0 net8 A0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN5 Y B0 net8 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMP3 net033 A0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MPM1 Y B0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MPM0 Y A1 net033 VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI21X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI21X6H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MNM1 net8 A1 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MNM0 net8 A0 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN5 Y B0 net8 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMP3 net033 A0 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MPM1 Y B0 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MPM0 Y A1 net033 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI21X8H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI21X8H7L A0 A1 B0 VDD VSS Y
*.PININFO A0:I A1:I B0:I Y:O VDD:B VSS:B
MNM1 net8 A1 VSS VSS nm1p2_lvt_lp W=1.2u L=60n m=1
MNM0 net8 A0 VSS VSS nm1p2_lvt_lp W=1.2u L=60n m=1
MMN5 Y B0 net8 VSS nm1p2_lvt_lp W=1.2u L=60n m=1
MMP3 net033 A0 VDD VDD pm1p2_lvt_lp W=1.52u L=60n m=1
MPM1 Y B0 VDD VDD pm1p2_lvt_lp W=1.52u L=60n m=1
MPM0 Y A1 net033 VDD pm1p2_lvt_lp W=1.52u L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI221X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI221X0P5H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MNM6 net31 B0 net39 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM5 net31 B1 net39 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM4 net39 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM7 Y C0 net31 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net39 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM4 Y B0 net22 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 Y A0 net18 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM7 Y C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM6 net18 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM5 net22 B1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI221X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI221X0P7H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MNM6 net31 B0 net39 VSS nm1p2_lvt_lp W=175n L=60n m=1
MNM5 net31 B1 net39 VSS nm1p2_lvt_lp W=175n L=60n m=1
MNM4 net39 A1 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MNM7 Y C0 net31 VSS nm1p2_lvt_lp W=175n L=60n m=1
MNM0 net39 A0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MPM4 Y B0 net22 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM1 Y A0 net18 VDD pm1p2_lvt_lp W=222n L=60n m=1
MPM7 Y C0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MPM6 net18 A1 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MPM5 net22 B1 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI221X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI221X1H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MNM6 net31 B0 net39 VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM5 net31 B1 net39 VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM4 net39 A1 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM7 Y C0 net31 VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM0 net39 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MPM4 Y B0 net22 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM1 Y A0 net18 VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM7 Y C0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM6 net18 A1 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM5 net22 B1 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI221X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI221X1P4H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MNM6 net31 B0 net39 VSS nm1p2_lvt_lp W=245n L=60n m=1
MNM5 net31 B1 net39 VSS nm1p2_lvt_lp W=245n L=60n m=1
MNM4 net39 A1 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MNM7 Y C0 net31 VSS nm1p2_lvt_lp W=245n L=60n m=1
MNM0 net39 A0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MPM4 Y B0 net22 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM1 Y A0 net18 VDD pm1p2_lvt_lp W=314n L=60n m=1
MPM7 Y C0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MPM6 net18 A1 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MPM5 net22 B1 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI221X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI221X2H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MNM6 net31 B0 net39 VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM5 net31 B1 net39 VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM4 net39 A1 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM7 Y C0 net31 VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM0 net39 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MPM4 Y B0 net22 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM1 Y A0 net18 VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM7 Y C0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM6 net18 A1 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM5 net22 B1 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI221X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI221X3H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MNM6 net31 B0 net39 VSS nm1p2_lvt_lp W=450n L=60n m=1
MNM5 net31 B1 net39 VSS nm1p2_lvt_lp W=450n L=60n m=1
MNM4 net39 A1 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MNM7 Y C0 net31 VSS nm1p2_lvt_lp W=450n L=60n m=1
MNM0 net39 A0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MPM4 Y B0 net22 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM1 Y A0 net18 VDD pm1p2_lvt_lp W=570n L=60n m=1
MPM7 Y C0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MPM6 net18 A1 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MPM5 net22 B1 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI221X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI221X4H7L A0 A1 B0 B1 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I Y:O VDD:B VSS:B
MNM6 net31 B0 net39 VSS nm1p2_lvt_lp W=600n L=60n m=1
MNM5 net31 B1 net39 VSS nm1p2_lvt_lp W=600n L=60n m=1
MNM4 net39 A1 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MNM7 Y C0 net31 VSS nm1p2_lvt_lp W=600n L=60n m=1
MNM0 net39 A0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MPM4 Y B0 net22 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM1 Y A0 net18 VDD pm1p2_lvt_lp W=760n L=60n m=1
MPM7 Y C0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MPM6 net18 A1 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MPM5 net22 B1 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI222X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI222X0P5H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 Y C1 net44 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM4 Y C0 net44 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 net44 B1 net52 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net44 B0 net52 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net52 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net52 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM5 Y C1 net11 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM4 net11 C0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 Y B1 net19 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net19 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 Y A1 net27 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net27 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI222X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI222X0P7H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 Y C1 net44 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM4 Y C0 net44 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM3 net44 B1 net52 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM2 net44 B0 net52 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM1 net52 A1 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM0 net52 A0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMPM5 Y C1 net11 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM4 net11 C0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM3 Y B1 net19 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM2 net19 B0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM1 Y A1 net27 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM0 net27 A0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI222X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI222X1H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 Y C1 net44 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM4 Y C0 net44 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM3 net44 B1 net52 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM2 net44 B0 net52 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM1 net52 A1 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM0 net52 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMPM5 Y C1 net11 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM4 net11 C0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM3 Y B1 net19 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM2 net19 B0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM1 Y A1 net27 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM0 net27 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI222X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI222X1P4H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 Y C1 net44 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM4 Y C0 net44 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM3 net44 B1 net52 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM2 net44 B0 net52 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM1 net52 A1 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM0 net52 A0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMPM5 Y C1 net11 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM4 net11 C0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM3 Y B1 net19 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM2 net19 B0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM1 Y A1 net27 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM0 net27 A0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI222X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI222X2H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 Y C1 net44 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM4 Y C0 net44 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM3 net44 B1 net52 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM2 net44 B0 net52 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM1 net52 A1 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM0 net52 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMPM5 Y C1 net11 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM4 net11 C0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM3 Y B1 net19 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM2 net19 B0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM1 Y A1 net27 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM0 net27 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI222X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI222X3H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 Y C1 net44 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM4 Y C0 net44 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM3 net44 B1 net52 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM2 net44 B0 net52 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM1 net52 A1 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM0 net52 A0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMPM5 Y C1 net11 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM4 net11 C0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM3 Y B1 net19 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM2 net19 B0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM1 Y A1 net27 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM0 net27 A0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI222X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI222X4H7L A0 A1 B0 B1 C0 C1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Y:O VDD:B VSS:B
MMNM5 Y C1 net44 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM4 Y C0 net44 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM3 net44 B1 net52 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM2 net44 B0 net52 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM1 net52 A1 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM0 net52 A0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMPM5 Y C1 net11 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM4 net11 C0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM3 Y B1 net19 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM2 net19 B0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM1 Y A1 net27 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM0 net27 A0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI22X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI22X0P5H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MNM0 Y B1 net8 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 net8 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net8 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 Y B0 net8 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP5 Y A1 net046 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM2 net046 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 Y B1 net049 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 net049 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI22X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI22X0P7H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MNM0 Y B1 net8 VSS nm1p2_lvt_lp W=175n L=60n m=1
MNM2 net8 A0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MNM1 net8 A1 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN5 Y B0 net8 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMP5 Y A1 net046 VDD pm1p2_lvt_lp W=222n L=60n m=1
MPM2 net046 A0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MPM0 Y B1 net049 VDD pm1p2_lvt_lp W=222n L=60n m=1
MPM1 net049 B0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI22X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI22X1H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MNM4 net8 A1 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM3 net8 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN5 Y B0 net8 VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM5 Y B1 net8 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMP5 Y A1 net046 VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM3 net046 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM5 Y B1 net049 VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM4 net049 B0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI22X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI22X1P4H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MNM0 Y B1 net8 VSS nm1p2_lvt_lp W=245n L=60n m=1
MNM2 net8 A0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MNM1 net8 A1 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN5 Y B0 net8 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMP5 Y A1 net046 VDD pm1p2_lvt_lp W=314n L=60n m=1
MPM2 net046 A0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MPM0 Y B1 net049 VDD pm1p2_lvt_lp W=314n L=60n m=1
MPM1 net049 B0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI22X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI22X2H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MNM3 net8 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM5 Y B1 net8 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN5 Y B0 net8 VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM4 net8 A1 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MPM4 Y B1 net049 VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM3 Y A1 net046 VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM5 net049 B0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM2 net046 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI22X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI22X3H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MNM3 net8 A0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MNM4 net8 A1 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MNM5 Y B1 net8 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMN5 Y B0 net8 VSS nm1p2_lvt_lp W=450n L=60n m=1
MPM4 Y B1 net049 VDD pm1p2_lvt_lp W=570n L=60n m=1
MPM5 net049 B0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MPM2 net046 A0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MPM3 Y A1 net046 VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI22X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI22X4H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MNM3 net8 A0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MNM4 net8 A1 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MNM5 Y B1 net8 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN5 Y B0 net8 VSS nm1p2_lvt_lp W=600n L=60n m=1
MPM4 Y B1 net049 VDD pm1p2_lvt_lp W=760n L=60n m=1
MPM5 net049 B0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MPM2 net046 A0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MPM3 Y A1 net046 VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI22X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI22X6H7L A0 A1 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I B0:I B1:I Y:O VDD:B VSS:B
MNM3 net8 A0 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MNM4 net8 A1 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MNM5 Y B1 net8 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN5 Y B0 net8 VSS nm1p2_lvt_lp W=900n L=60n m=1
MPM4 Y B1 net049 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MPM5 net049 B0 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MPM2 net046 A0 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MPM3 Y A1 net046 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2BB1X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2BB1X0P5H7L A0N A1N B0 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I Y:O VDD:B VSS:B
MMN7 net042 A1N net45 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net45 A0N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 Y net042 net42 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 net42 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP7 net042 A0N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net042 A1N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 Y net042 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM2 Y B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2BB1X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2BB1X0P7H7L A0N A1N B0 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I Y:O VDD:B VSS:B
MMN7 net042 A1N net45 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net45 A0N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 Y net042 net42 VSS nm1p2_lvt_lp W=175n L=60n m=1
MNM2 net42 B0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMP7 net042 A0N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net042 A1N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 Y net042 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MPM2 Y B0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2BB1X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2BB1X1H7L A0N A1N B0 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I Y:O VDD:B VSS:B
MMN7 net042 A1N net45 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net42 B0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM0 net45 A0N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN10 Y net042 net42 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMP7 net042 A0N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net042 A1N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP9 Y net042 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM1 Y B0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2BB1X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2BB1X1P4H7L A0N A1N B0 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I Y:O VDD:B VSS:B
MMN7 net042 A1N net45 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net45 A0N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 Y net042 net42 VSS nm1p2_lvt_lp W=245n L=60n m=1
MNM2 net42 B0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMP7 net042 A0N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net042 A1N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 Y net042 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MPM2 Y B0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2BB1X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2BB1X2H7L A0N A1N B0 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I Y:O VDD:B VSS:B
MMN7 net042 A1N net45 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net42 B0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM0 net45 A0N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN10 Y net042 net42 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP9 Y net042 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP5 net042 A1N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 Y B0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM0 net042 A0N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2BB1X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2BB1X3H7L A0N A1N B0 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I Y:O VDD:B VSS:B
MMN7 net042 A1N net45 VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM2 net45 A0N VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM1 net42 B0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MNM0 Y net042 net42 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMP9 Y net042 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP5 net042 A1N VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM1 Y B0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MPM0 net042 A0N VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2BB1X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2BB1X4H7L A0N A1N B0 VDD VSS Z
*.PININFO A0N:I A1N:I B0:I Z:O VDD:B VSS:B
MMN7 net042 A1N net45 VSS nm1p2_lvt_lp W=250n L=60n m=1
MNM2 net45 A0N VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MNM1 net42 B0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MNM0 Z net042 net42 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMP9 Z net042 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP5 net042 A1N VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MPM1 Z B0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MPM0 net042 A0N VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2BB1X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2BB1X6H7L A0N A1N B0 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I Y:O VDD:B VSS:B
MMN7 net042 A1N net45 VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM2 net45 A0N VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM1 net42 B0 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MNM0 Y net042 net42 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMP9 Y net042 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP5 net042 A1N VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM1 Y B0 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MPM0 net042 A0N VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2BB2X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2BB2X0P5H7L A0N A1N B0 B1 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I B1:I Y:O VDD:B VSS:B
MNM3 net8 B1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 Y net35 net8 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net8 B0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net48 A1N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN10 net35 A0N net48 VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM2 net058 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 Y net35 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP8 net35 A0N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM3 Y B1 net058 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net35 A1N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2BB2X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2BB2X0P7H7L A0N A1N B0 B1 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I B1:I Y:O VDD:B VSS:B
MNM3 net8 B1 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MNM2 Y net35 net8 VSS nm1p2_lvt_lp W=175n L=60n m=1
MNM1 net8 B0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MNM0 net48 A1N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN10 net35 A0N net48 VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM2 net058 B0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MPM1 Y net35 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMP8 net35 A0N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM3 Y B1 net058 VDD pm1p2_lvt_lp W=222n L=60n m=1
MPM0 net35 A1N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2BB2X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2BB2X1H7L A0N A1N B0 B1 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I B1:I Y:O VDD:B VSS:B
MNM5 net8 B1 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM2 Y net35 net8 VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM4 net8 B0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM0 net48 A1N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN10 net35 A0N net48 VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM5 Y B1 net058 VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM1 Y net35 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP8 net35 A0N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM4 net058 B0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM0 net35 A1N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2BB2X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2BB2X1P4H7L A0N A1N B0 B1 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I B1:I Y:O VDD:B VSS:B
MNM3 net8 B1 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MNM2 Y net35 net8 VSS nm1p2_lvt_lp W=245n L=60n m=1
MNM1 net8 B0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MNM0 net48 A1N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN10 net35 A0N net48 VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM2 net058 B0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MPM1 Y net35 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMP8 net35 A0N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM3 Y B1 net058 VDD pm1p2_lvt_lp W=314n L=60n m=1
MPM0 net35 A1N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2BB2X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2BB2X2H7L A0N A1N B0 B1 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I B1:I Y:O VDD:B VSS:B
MNM4 net8 B0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM2 Y net35 net8 VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM5 net8 B1 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM0 net48 A1N VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN10 net35 A0N net48 VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM5 Y B1 net058 VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM1 Y net35 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP8 net35 A0N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM4 net058 B0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM0 net35 A1N VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2BB2X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2BB2X3H7L A0N A1N B0 B1 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I B1:I Y:O VDD:B VSS:B
MNM6 net8 B1 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MNM5 net8 B0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MNM2 Y net35 net8 VSS nm1p2_lvt_lp W=450n L=60n m=1
MNM4 net48 A1N VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN10 net35 A0N net48 VSS nm1p2_lvt_lp W=210n L=60n m=1
MPM6 Y B1 net058 VDD pm1p2_lvt_lp W=570n L=60n m=1
MPM1 Y net35 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMP8 net35 A0N VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM5 net058 B0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MPM4 net35 A1N VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2BB2X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2BB2X4H7L A0N A1N B0 B1 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I B1:I Y:O VDD:B VSS:B
MNM6 net8 B1 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MNM5 net8 B0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MNM2 Y net35 net8 VSS nm1p2_lvt_lp W=600n L=60n m=1
MNM4 net48 A1N VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMN10 net35 A0N net48 VSS nm1p2_lvt_lp W=250n L=60n m=1
MPM6 Y B1 net058 VDD pm1p2_lvt_lp W=760n L=60n m=1
MPM1 Y net35 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP8 net35 A0N VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MPM5 net058 B0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MPM4 net35 A1N VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2BB2X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2BB2X6H7L A0N A1N B0 B1 VDD VSS Y
*.PININFO A0N:I A1N:I B0:I B1:I Y:O VDD:B VSS:B
MNM6 net8 B1 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MNM5 net8 B0 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MNM2 Y net35 net8 VSS nm1p2_lvt_lp W=900n L=60n m=1
MNM4 net48 A1N VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN10 net35 A0N net48 VSS nm1p2_lvt_lp W=300n L=60n m=1
MPM6 Y B1 net058 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MPM1 Y net35 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP8 net35 A0N VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM5 net058 B0 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MPM4 net35 A1N VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2XB1X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2XB1X0P5H7L A0 A1N B0 VDD VSS Y
*.PININFO A0:I A1N:I B0:I Y:O VDD:B VSS:B
MMNM2 Y B0 net17 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net17 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net17 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM1 Y A1 net12 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 Y B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net12 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 A1N VDD VSS A1 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2XB1X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2XB1X0P7H7L A0 A1N B0 VDD VSS Y
*.PININFO A0:I A1N:I B0:I Y:O VDD:B VSS:B
MMNM2 Y B0 net17 VSS nm1p2_lvt_lp W=174n L=60n m=1
MMNM1 net17 A1 VSS VSS nm1p2_lvt_lp W=174n L=60n m=1
MMNM0 net17 A0 VSS VSS nm1p2_lvt_lp W=174n L=60n m=1
MMPM1 Y A1 net12 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM2 Y B0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM0 net12 A0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
XXI3 A1N VDD VSS A1 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2XB1X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2XB1X1H7L A0 A1N B0 VDD VSS Y
*.PININFO A0:I A1N:I B0:I Y:O VDD:B VSS:B
MMNM2 Y B0 net17 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM1 net17 A1 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM0 net17 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMPM1 Y A1 net12 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM2 Y B0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM0 net12 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
XXI3 A1N VDD VSS A1 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2XB1X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2XB1X1P4H7L A0 A1N B0 VDD VSS Y
*.PININFO A0:I A1N:I B0:I Y:O VDD:B VSS:B
MMNM2 Y B0 net17 VSS nm1p2_lvt_lp W=246n L=60n m=1
MMNM1 net17 A1 VSS VSS nm1p2_lvt_lp W=246n L=60n m=1
MMNM0 net17 A0 VSS VSS nm1p2_lvt_lp W=246n L=60n m=1
MMPM1 Y A1 net12 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM2 Y B0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM0 net12 A0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
XXI3 A1N VDD VSS A1 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2XB1X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2XB1X2H7L A0 A1N B0 VDD VSS Y
*.PININFO A0:I A1N:I B0:I Y:O VDD:B VSS:B
MMNM2 Y B0 net17 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM1 net17 A1 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM0 net17 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMPM1 Y A1 net12 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM2 Y B0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM0 net12 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
XXI3 A1N VDD VSS A1 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2XB1X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2XB1X3H7L A0 A1N B0 VDD VSS Y
*.PININFO A0:I A1N:I B0:I Y:O VDD:B VSS:B
MMNM2 Y B0 net17 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM1 net17 A1 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM0 net17 A0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMPM1 Y A1 net12 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM2 Y B0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM0 net12 A0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
XXI3 A1N VDD VSS A1 / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2XB1X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2XB1X4H7L A0 A1N B0 VDD VSS Y
*.PININFO A0:I A1N:I B0:I Y:O VDD:B VSS:B
MMNM2 Y B0 net17 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM1 net17 A1 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM0 net17 A0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMPM1 Y A1 net12 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM2 Y B0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM0 net12 A0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
XXI3 A1N VDD VSS A1 / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI2XB1X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI2XB1X6H7L A0 A1N B0 VDD VSS Y
*.PININFO A0:I A1N:I B0:I Y:O VDD:B VSS:B
MMNM2 Y B0 net17 VSS nm1p2_lvt_lp W=900n L=60n m=1
MMNM1 net17 A1 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMNM0 net17 A0 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMPM1 Y A1 net12 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMPM2 Y B0 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMPM0 net12 A0 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
XXI3 A1N VDD VSS A1 / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI31X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI31X0P5H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMNM3 Y B0 net34 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net34 A2 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net34 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net34 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM2 net17 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 Y B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 net13 A1 net17 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 Y A2 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI31X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI31X0P7H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMNM3 Y B0 net34 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM2 net34 A2 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM1 net34 A1 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM0 net34 A0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MPM2 net17 A0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM3 Y B0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MPM1 net13 A1 net17 VDD pm1p2_lvt_lp W=222n L=60n m=1
MPM0 Y A2 net13 VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI31X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI31X1H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMNM3 Y B0 net34 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM2 net34 A2 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM1 net34 A1 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM0 net34 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MPM2 net17 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM3 Y B0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM1 net13 A1 net17 VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM0 Y A2 net13 VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI31X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI31X1P4H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMNM3 Y B0 net34 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM2 net34 A2 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM1 net34 A1 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM0 net34 A0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MPM2 net17 A0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM3 Y B0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MPM1 net13 A1 net17 VDD pm1p2_lvt_lp W=314n L=60n m=1
MPM0 Y A2 net13 VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI31X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI31X2H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMNM3 Y B0 net34 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM2 net34 A2 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM1 net34 A1 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM0 net34 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MPM2 net17 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM3 Y B0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM1 net13 A1 net17 VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM0 Y A2 net13 VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI31X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI31X3H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMNM3 Y B0 net34 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM2 net34 A2 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM1 net34 A1 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM0 net34 A0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MPM2 net17 A0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM3 Y B0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MPM1 net13 A1 net17 VDD pm1p2_lvt_lp W=570n L=60n m=1
MPM0 Y A2 net13 VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI31X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI31X4H7L A0 A1 A2 B0 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I Y:O VDD:B VSS:B
MMNM3 Y B0 net34 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM2 net34 A2 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM1 net34 A1 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM0 net34 A0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MPM2 net17 A0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM3 Y B0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MPM1 net13 A1 net17 VDD pm1p2_lvt_lp W=760n L=60n m=1
MPM0 Y A2 net13 VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI32X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI32X0P5H7L A0 A1 A2 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I Y:O VDD:B VSS:B
MMNM4 Y B1 net42 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 Y B0 net42 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net42 A2 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net42 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net42 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM4 Y B1 net21 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net21 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 Y A2 net9 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net9 A1 net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI32X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI32X0P7H7L A0 A1 A2 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I Y:O VDD:B VSS:B
MMNM4 Y B1 net42 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM3 Y B0 net42 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM2 net42 A2 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM1 net42 A1 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM0 net42 A0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMPM4 Y B1 net21 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM3 net21 B0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM2 Y A2 net9 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM1 net9 A1 net13 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI32X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI32X1H7L A0 A1 A2 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I Y:O VDD:B VSS:B
MMNM4 Y B1 net42 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM3 Y B0 net42 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM2 net42 A2 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM1 net42 A1 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM0 net42 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMPM4 Y B1 net21 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM3 net21 B0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM2 Y A2 net9 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM1 net9 A1 net13 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI32X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI32X1P4H7L A0 A1 A2 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I Y:O VDD:B VSS:B
MMNM4 Y B1 net42 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM3 Y B0 net42 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM2 net42 A2 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM1 net42 A1 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM0 net42 A0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMPM4 Y B1 net21 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM3 net21 B0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM2 Y A2 net9 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM1 net9 A1 net13 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI32X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI32X2H7L A0 A1 A2 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I Y:O VDD:B VSS:B
MMNM4 Y B1 net42 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM3 Y B0 net42 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM2 net42 A2 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM1 net42 A1 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM0 net42 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMPM4 Y B1 net21 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM3 net21 B0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM2 Y A2 net9 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM1 net9 A1 net13 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI32X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI32X3H7L A0 A1 A2 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I Y:O VDD:B VSS:B
MMNM4 Y B1 net42 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM3 Y B0 net42 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM2 net42 A2 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM1 net42 A1 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM0 net42 A0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMPM4 Y B1 net21 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM3 net21 B0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM2 Y A2 net9 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM1 net9 A1 net13 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI32X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI32X4H7L A0 A1 A2 B0 B1 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I Y:O VDD:B VSS:B
MMNM4 Y B1 net42 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM3 Y B0 net42 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM2 net42 A2 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM1 net42 A1 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM0 net42 A0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMPM4 Y B1 net21 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM3 net21 B0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM2 Y A2 net9 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM1 net9 A1 net13 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM0 net13 A0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI33X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI33X0P5H7L A0 A1 A2 B0 B1 B2 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I B2:I Y:O VDD:B VSS:B
MMNM5 Y B2 net52 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM4 Y B1 net52 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM3 Y B0 net52 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM2 net52 A2 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM1 net52 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net52 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM5 Y B2 net15 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM4 net15 B1 net23 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM3 net23 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 Y A2 net11 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net11 A1 net19 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net19 A0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI33X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI33X0P7H7L A0 A1 A2 B0 B1 B2 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I B2:I Y:O VDD:B VSS:B
MMNM5 Y B2 net52 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM4 Y B1 net52 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM3 Y B0 net52 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM2 net52 A2 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM1 net52 A1 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMNM0 net52 A0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMPM5 Y B2 net15 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM4 net15 B1 net23 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM3 net23 B0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM2 Y A2 net11 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM1 net11 A1 net19 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM0 net19 A0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI33X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI33X1H7L A0 A1 A2 B0 B1 B2 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I B2:I Y:O VDD:B VSS:B
MMNM5 Y B2 net52 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM4 Y B1 net52 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM3 Y B0 net52 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM2 net52 A2 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM1 net52 A1 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM0 net52 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMPM5 Y B2 net15 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM4 net15 B1 net23 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM3 net23 B0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM2 Y A2 net11 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM1 net11 A1 net19 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM0 net19 A0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI33X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI33X1P4H7L A0 A1 A2 B0 B1 B2 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I B2:I Y:O VDD:B VSS:B
MMNM5 Y B2 net52 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM4 Y B1 net52 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM3 Y B0 net52 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM2 net52 A2 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM1 net52 A1 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMNM0 net52 A0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMPM5 Y B2 net15 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM4 net15 B1 net23 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM3 net23 B0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM2 Y A2 net11 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM1 net11 A1 net19 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM0 net19 A0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI33X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI33X2H7L A0 A1 A2 B0 B1 B2 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I B2:I Y:O VDD:B VSS:B
MMNM5 Y B2 net52 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM4 Y B1 net52 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM3 Y B0 net52 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM2 net52 A2 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM1 net52 A1 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM0 net52 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMPM5 Y B2 net15 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM4 net15 B1 net23 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM3 net23 B0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM2 Y A2 net11 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM1 net11 A1 net19 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM0 net19 A0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI33X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI33X3H7L A0 A1 A2 B0 B1 B2 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I B2:I Y:O VDD:B VSS:B
MMNM5 Y B2 net52 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM4 Y B1 net52 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM3 Y B0 net52 VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM2 net52 A2 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM1 net52 A1 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMNM0 net52 A0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMPM5 Y B2 net15 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM4 net15 B1 net23 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM3 net23 B0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM2 Y A2 net11 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM1 net11 A1 net19 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMPM0 net19 A0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAI33X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAI33X4H7L A0 A1 A2 B0 B1 B2 VDD VSS Y
*.PININFO A0:I A1:I A2:I B0:I B1:I B2:I Y:O VDD:B VSS:B
MMNM5 Y B2 net52 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM4 Y B1 net52 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM3 Y B0 net52 VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM2 net52 A2 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM1 net52 A1 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMNM0 net52 A0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMPM5 Y B2 net15 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM4 net15 B1 net23 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM3 net23 B0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM2 Y A2 net11 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM1 net11 A1 net19 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMPM0 net19 A0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAO211X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAO211X0P5H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM6 net26 C0 net14 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM5 net14 A0 net17 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM0 net17 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM4 net14 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM7 net26 C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM3 net34 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM2 net34 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM8 net26 B0 net34 VSS nm1p2_lvt_lp W=150n L=60n m=1
XXI3 net26 VDD VSS Y / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAO211X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAO211X0P7H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM6 net26 C0 net14 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM5 net14 A0 net17 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM0 net17 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM4 net14 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM7 net26 C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM3 net34 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM2 net34 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM8 net26 B0 net34 VSS nm1p2_lvt_lp W=150n L=60n m=1
XXI3 net26 VDD VSS Y / INV pl=6e-08 pw=2.22e-07 nl=6e-08 nw=1.74e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAO211X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAO211X1H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM6 net26 C0 net14 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM5 net14 A0 net17 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM0 net17 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM4 net14 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM7 net26 C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM3 net34 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM2 net34 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM8 net26 B0 net34 VSS nm1p2_lvt_lp W=150n L=60n m=1
XXI3 net26 VDD VSS Y / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAO211X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAO211X1P4H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM6 net26 C0 net14 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM5 net14 A0 net17 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM0 net17 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM4 net14 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM7 net26 C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM3 net34 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM2 net34 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM8 net26 B0 net34 VSS nm1p2_lvt_lp W=150n L=60n m=1
XXI3 net26 VDD VSS Y / INV pl=6e-08 pw=3.14e-07 nl=6e-08 nw=2.46e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAO211X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAO211X2H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM6 net26 C0 net14 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM5 net14 A0 net17 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM0 net17 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM4 net14 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM7 net26 C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM3 net34 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM2 net34 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM8 net26 B0 net34 VSS nm1p2_lvt_lp W=150n L=60n m=1
XXI0 net26 VDD VSS Y / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAO211X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAO211X3H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM6 net26 C0 net14 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMM5 net14 A0 net17 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMM0 net17 A1 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMM4 net14 B0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMM7 net26 C0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMM3 net34 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMM2 net34 A1 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMM8 net26 B0 net34 VSS nm1p2_lvt_lp W=210n L=60n m=1
XXI3 net26 VDD VSS Y / INV pl=6e-08 pw=5.7e-07 nl=6e-08 nw=4.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAO211X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAO211X4H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM6 net26 C0 net14 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMM5 net14 A0 net17 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMM0 net17 A1 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MMM4 net14 B0 VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MMM7 net26 C0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMM3 net34 A0 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMM2 net34 A1 VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMM8 net26 B0 net34 VSS nm1p2_lvt_lp W=250n L=60n m=1
XXI3 net26 VDD VSS Y / INV pl=6e-08 pw=7.6e-07 nl=6e-08 nw=6e-07
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAOI211X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAOI211X0P5H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM7 Y C0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM3 net10 A0 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM2 net10 A1 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMM8 Y B0 net10 VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM0 Y C0 net26 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM5 net26 A0 net29 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM0 net29 A1 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
MMM4 net26 B0 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAOI211X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAOI211X0P7H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM7 Y C0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMM3 net10 A0 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMM2 net10 A1 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMM8 Y B0 net10 VSS nm1p2_lvt_lp W=175n L=60n m=1
MPM0 Y C0 net26 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMM5 net26 A0 net29 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMM0 net29 A1 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
MMM4 net26 B0 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAOI211X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAOI211X1H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM7 Y C0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMM3 net10 A0 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMM2 net10 A1 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMM8 Y B0 net10 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMM6 Y C0 net26 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMM5 net26 A0 net29 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMM0 net29 A1 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MMM4 net26 B0 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAOI211X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAOI211X1P4H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM7 Y C0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMM3 net10 A0 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMM2 net10 A1 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMM8 Y B0 net10 VSS nm1p2_lvt_lp W=245n L=60n m=1
MPM0 Y C0 net26 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMM5 net26 A0 net29 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMM0 net29 A1 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
MMM4 net26 B0 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAOI211X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAOI211X2H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM7 Y C0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMM3 net10 A0 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMM2 net10 A1 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMM8 Y B0 net10 VSS nm1p2_lvt_lp W=300n L=60n m=1
MPM0 Y C0 net26 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMM5 net26 A0 net29 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMM0 net29 A1 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMM4 net26 B0 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAOI211X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAOI211X3H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM7 Y C0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMM3 net10 A0 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMM2 net10 A1 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MMM8 Y B0 net10 VSS nm1p2_lvt_lp W=450n L=60n m=1
MPM0 Y C0 net26 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMM5 net26 A0 net29 VDD pm1p2_lvt_lp W=570n L=60n m=1
MMM0 net29 A1 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MMM4 net26 B0 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OAOI211X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OAOI211X4H7L A0 A1 B0 C0 VDD VSS Y
*.PININFO A0:I A1:I B0:I C0:I Y:O VDD:B VSS:B
MMM7 Y C0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMM3 net10 A0 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMM2 net10 A1 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMM8 Y B0 net10 VSS nm1p2_lvt_lp W=600n L=60n m=1
MPM0 Y C0 net26 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMM5 net26 A0 net29 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMM0 net29 A1 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MMM4 net26 B0 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR2X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR2X0P5H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN2 net21 B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 net21 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP2 net21 B net016 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 net016 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI4 net21 VDD VSS Y / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR2X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR2X0P7H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN2 net21 B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 net21 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP2 net21 B net016 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 net016 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI4 net21 VDD VSS Y / INV pl=6e-08 pw=2.22e-07 nl=6e-08 nw=1.74e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR2X12H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR2X12H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN2 net21 B VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMN0 net21 A VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MMP2 net21 B net016 VDD pm1p2_lvt_lp W=760n L=60n m=1
MMP1 net016 A VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
XXI4 net21 VDD VSS Y / INV pl=6e-08 pw=22.8e-07 nl=6e-08 nw=18e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR2X16H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR2X16H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN2 net21 B VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMN0 net21 A VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MMP2 net21 B net016 VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MMP1 net016 A VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
XXI4 net21 VDD VSS Y / INV pl=6e-08 pw=30.4e-07 nl=6e-08 nw=24e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR2X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR2X1H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN2 net21 B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 net21 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP2 net21 B net016 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 net016 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI4 net21 VDD VSS Y / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR2X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR2X1P4H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN2 net21 B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 net21 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP2 net21 B net016 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 net016 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI4 net21 VDD VSS Y / INV pl=6e-08 pw=3.14e-07 nl=6e-08 nw=2.46e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR2X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR2X2H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN2 net21 B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 net21 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP2 net21 B net016 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMP1 net016 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI4 net21 VDD VSS Y / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR2X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR2X3H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN2 net21 B VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN0 net21 A VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMP2 net21 B net016 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMP1 net016 A VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
XXI4 net21 VDD VSS Y / INV pl=6e-08 pw=5.7e-07 nl=6e-08 nw=4.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR2X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR2X4H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN2 net21 B VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMN0 net21 A VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMP2 net21 B net016 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMP1 net016 A VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
XXI4 net21 VDD VSS Y / INV pl=6e-08 pw=7.6e-07 nl=6e-08 nw=6e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR2X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR2X6H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN2 net21 B VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN0 net21 A VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP2 net21 B net016 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMP1 net016 A VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
XXI4 net21 VDD VSS Y / INV pl=6e-08 pw=11.4e-07 nl=6e-08 nw=9e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR2X8H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR2X8H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN2 net21 B VSS VSS nm1p2_lvt_lp W=500n L=60n m=1
MMN0 net21 A VSS VSS nm1p2_lvt_lp W=500n L=60n m=1
MMP2 net21 B net016 VDD pm1p2_lvt_lp W=620n L=60n m=1
MMP1 net016 A VDD VDD pm1p2_lvt_lp W=620n L=60n m=1
XXI4 net21 VDD VSS Y / INV pl=6e-08 pw=15.2e-07 nl=6e-08 nw=12e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR3X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR3X0P5H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MNM0 net27 B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net27 C VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN3 net27 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP3 net27 C net22 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net22 B net020 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 net020 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI4 net27 VDD VSS Y / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR3X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR3X0P7H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MNM0 net27 B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net27 C VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN3 net27 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP3 net27 C net22 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net22 B net020 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 net020 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI4 net27 VDD VSS Y / INV pl=6e-08 pw=2.22e-07 nl=6e-08 nw=1.74e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR3X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR3X1H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MNM0 net27 B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net27 C VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN3 net27 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP3 net27 C net22 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net22 B net020 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 net020 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI4 net27 VDD VSS Y / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR3X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR3X1P4H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MNM0 net27 B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net27 C VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN3 net27 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP3 net27 C net22 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net22 B net020 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 net020 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI4 net27 VDD VSS Y / INV pl=6e-08 pw=3.14e-07 nl=6e-08 nw=2.46e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR3X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR3X2H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MNM0 net27 B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net27 C VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN3 net27 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP3 net27 C net22 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM0 net22 B net020 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 net020 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI4 net27 VDD VSS Y / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR3X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR3X3H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MNM0 net27 B VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM1 net27 C VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN3 net27 A VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMP3 net27 C net22 VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM0 net22 B net020 VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM1 net020 A VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
XXI4 net27 VDD VSS Y / INV pl=6e-08 pw=5.7e-07 nl=6e-08 nw=4.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR3X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR3X4H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MNM0 net27 B VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MNM1 net27 C VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMN3 net27 A VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMP3 net27 C net22 VDD pm1p2_lvt_lp W=310n L=60n m=1
MPM0 net22 B net020 VDD pm1p2_lvt_lp W=310n L=60n m=1
MPM1 net020 A VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
XXI4 net27 VDD VSS Y / INV pl=6e-08 pw=7.6e-07 nl=6e-08 nw=6e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR3X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR3X6H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MNM0 net27 B VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM1 net27 C VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN3 net27 A VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMP3 net27 C net22 VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM0 net22 B net020 VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM1 net020 A VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
XXI4 net27 VDD VSS Y / INV pl=6e-08 pw=11.4e-07 nl=6e-08 nw=9e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR3X8H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR3X8H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MNM0 net27 B VSS VSS nm1p2_lvt_lp W=500n L=60n m=1
MNM1 net27 C VSS VSS nm1p2_lvt_lp W=500n L=60n m=1
MMN3 net27 A VSS VSS nm1p2_lvt_lp W=500n L=60n m=1
MMP3 net27 C net22 VDD pm1p2_lvt_lp W=620n L=60n m=1
MPM0 net22 B net020 VDD pm1p2_lvt_lp W=620n L=60n m=1
MPM1 net020 A VDD VDD pm1p2_lvt_lp W=620n L=60n m=1
XXI4 net27 VDD VSS Y / INV pl=6e-08 pw=15.2e-07 nl=6e-08 nw=12e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR4X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR4X0P5H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MNM0 net22 B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net22 C VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 net22 D VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net22 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM3 net22 D net21 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net21 C net17 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net17 B net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net13 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI4 net22 VDD VSS Y / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR4X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR4X0P7H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MNM0 net22 B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net22 C VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 net22 D VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net22 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM3 net22 D net21 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net21 C net17 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net17 B net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net13 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI4 net22 VDD VSS Y / INV pl=6e-08 pw=2.22e-07 nl=6e-08 nw=1.74e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR4X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR4X1H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MNM0 net22 B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net22 C VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 net22 D VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net22 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM3 net22 D net21 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net21 C net17 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net17 B net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net13 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI4 net22 VDD VSS Y / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR4X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR4X1P4H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MNM0 net22 B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net22 C VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 net22 D VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net22 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM3 net22 D net21 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net21 C net17 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net17 B net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net13 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI4 net22 VDD VSS Y / INV pl=6e-08 pw=3.14e-07 nl=6e-08 nw=2.46e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR4X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR4X2H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MNM0 net22 B VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net22 C VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 net22 D VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMNM0 net22 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM3 net22 D net21 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM2 net21 C net17 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM1 net17 B net13 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net13 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI4 net22 VDD VSS Y / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR4X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR4X3H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MNM0 net22 B VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM1 net22 C VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM2 net22 D VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMNM0 net22 A VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMPM3 net22 D net21 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM2 net21 C net17 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM1 net17 B net13 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM0 net13 A VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
XXI4 net22 VDD VSS Y / INV pl=6e-08 pw=5.7e-07 nl=6e-08 nw=4.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR4X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR4X4H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MNM0 net22 B VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MNM1 net22 C VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MNM2 net22 D VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMNM0 net22 A VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMPM3 net22 D net21 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM2 net21 C net17 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM1 net17 B net13 VDD pm1p2_lvt_lp W=310n L=60n m=1
MMPM0 net13 A VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
XXI4 net22 VDD VSS Y / INV pl=6e-08 pw=7.6e-07 nl=6e-08 nw=6e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    OR4X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT OR4X6H7L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MNM0 net22 B VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM1 net22 C VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM2 net22 D VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMNM0 net22 A VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMPM3 net22 D net21 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM2 net21 C net17 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM1 net17 B net13 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM0 net13 A VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
XXI4 net22 VDD VSS Y / INV pl=6e-08 pw=11.4e-07 nl=6e-08 nw=9e-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFNQX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFNQX1H7L CKN D Q SE SI VDD VSS
*.PININFO CKN:I D:I SE:I SI:I Q:O VDD:B VSS:B
XXI9 net44 c cn VDD VSS net51 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI21 D SEN SE VDD VSS net76 / TSINV pl=60n pw=200n nl=60n nw=160n
XXI22 SI SE SEN VDD VSS net76 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI15 net48 cn c VDD VSS net51 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI14 net44 c cn VDD VSS net39 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI23 SE VDD VSS SEN / INV pl=60n pw=210n nl=60n nw=170n
XXI10 net51 VDD VSS net48 / INV pl=60n pw=190n nl=60n nw=150n
XXI12 net51 VDD VSS Q / INV pl=60n pw=270n nl=60n nw=210n
XXI4 CKN VDD VSS c / INV pl=60n pw=210n nl=60n nw=170n
XXI7 net39 VDD VSS net44 / INV pl=60n pw=190n nl=60n nw=150n
XXI13 c VDD VSS cn / INV pl=60n pw=210n nl=60n nw=170n
XXI6 cn c net76 net39 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFNQX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFNQX2H7L CKN D Q SE SI VDD VSS
*.PININFO CKN:I D:I SE:I SI:I Q:O VDD:B VSS:B
XXI14 net44 c cn VDD VSS net39 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI15 net48 cn c VDD VSS net51 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI22 SI SE SEN VDD VSS net76 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI21 D SEN SE VDD VSS net76 / TSINV pl=60n pw=210n nl=60n nw=170n
XXI9 net44 c cn VDD VSS net51 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI13 c VDD VSS cn / INV pl=60n pw=210n nl=60n nw=170n
XXI7 net39 VDD VSS net44 / INV pl=60n pw=200n nl=60n nw=160n
XXI4 CKN VDD VSS c / INV pl=60n pw=210n nl=60n nw=170n
XXI12 net51 VDD VSS Q / INV pl=60n pw=380n nl=60n nw=300n
XXI10 net51 VDD VSS net48 / INV pl=60n pw=210n nl=60n nw=170n
XXI23 SE VDD VSS SEN / INV pl=60n pw=210n nl=60n nw=170n
XXI6 cn c net76 net39 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFNQX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFNQX3H7L CKN D Q SE SI VDD VSS
*.PININFO CKN:I D:I SE:I SI:I Q:O VDD:B VSS:B
XXI13 c VDD VSS cn / INV pl=60n pw=210n nl=60n nw=170n
XXI10 net51 VDD VSS net48 / INV pl=60n pw=250n nl=60n nw=200n
XXI23 SE VDD VSS SEN / INV pl=60n pw=210n nl=60n nw=170n
XXI7 net39 VDD VSS net44 / INV pl=60n pw=210n nl=60n nw=170n
XXI4 CKN VDD VSS c / INV pl=60n pw=210n nl=60n nw=170n
XXI12 net51 VDD VSS Q / INV pl=60n pw=570n nl=60n nw=450n
XXI15 net48 cn c VDD VSS net51 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI9 net44 c cn VDD VSS net51 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI21 D SEN SE VDD VSS net76 / TSINV pl=60n pw=210n nl=60n nw=170n
XXI22 SI SE SEN VDD VSS net76 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI14 net44 c cn VDD VSS net39 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI6 cn c net76 net39 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFNRX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFNRX0P5H7L CKN D Q QN RN SE SI VDD VSS
*.PININFO CKN:I D:I RN:I SE:I SI:I Q:O QN:O VDD:B VSS:B
MMN1 net099 cn net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0147 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net099 r VSS VSS nm1p2_lvt_lp W=240n L=60n m=1
MMN4 net46 net33 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMP4 net54 r VDD VDD pm1p2_lvt_lp W=280n L=60n m=1
MMP2 net67 net0147 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net099 c net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=280n L=60n m=1
XXI29 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI33 SI SE SEN VDD VSS net076 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI30 D SEN SE VDD VSS net076 / TSINV pl=60n pw=280n nl=60n nw=240n
XXI9 c cn net46 net099 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
XXI32 cn c net076 net33 VDD VSS / TG pl=60n pw=260n nl=60n nw=200n
XXI34 SE VDD VSS SEN / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net099 VDD VSS QN / INV pl=60n pw=280n nl=60n nw=200n
XXI31 RN VDD VSS r / INV pl=60n pw=280n nl=60n nw=200n
XXI5 net0147 VDD VSS Q / INV pl=60n pw=280n nl=60n nw=200n
XXI13 c VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net099 VDD VSS net0147 / INV pl=60n pw=280n nl=60n nw=240n
XXI4 CKN VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFNRX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFNRX1H7L CKN D Q QN RN SE SI VDD VSS
*.PININFO CKN:I D:I RN:I SE:I SI:I Q:O QN:O VDD:B VSS:B
MNM2 net099 r VSS VSS nm1p2_lvt_lp W=240n L=60n m=1
MNM1 net53 net0147 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net099 cn net53 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 VSS VSS nm1p2_lvt_lp W=220n L=60n m=1
MPM2 net099 c net48 VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM1 net48 net0147 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM0 net54 r VDD VDD pm1p2_lvt_lp W=280n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=300n L=60n m=1
XXI29 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI33 SI SE SEN VDD VSS net076 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI30 D SEN SE VDD VSS net076 / TSINV pl=60n pw=280n nl=60n nw=240n
XXI9 c cn net46 net099 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
XXI32 cn c net076 net33 VDD VSS / TG pl=60n pw=260n nl=60n nw=200n
XXI34 SE VDD VSS SEN / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net099 VDD VSS QN / INV pl=60n pw=340n nl=60n nw=240n
XXI31 RN VDD VSS r / INV pl=60n pw=280n nl=60n nw=200n
XXI5 net0147 VDD VSS Q / INV pl=60n pw=340n nl=60n nw=240n
XXI13 c VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net099 VDD VSS net0147 / INV pl=60n pw=280n nl=60n nw=240n
XXI4 CKN VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFNRX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFNRX2H7L CKN D Q QN RN SE SI VDD VSS
*.PININFO CKN:I D:I RN:I SE:I SI:I Q:O QN:O VDD:B VSS:B
MMN1 net099 cn net66 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net66 net0147 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net099 r VSS VSS nm1p2_lvt_lp W=260n L=60n m=1
MMN4 net46 net33 VSS VSS nm1p2_lvt_lp W=240n L=60n m=1
MMP4 net54 r VDD VDD pm1p2_lvt_lp W=320n L=60n m=1
MMP2 net67 net0147 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net099 c net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=340n L=60n m=1
XXI29 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI33 SI SE SEN VDD VSS net076 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI30 D SEN SE VDD VSS net076 / TSINV pl=60n pw=280n nl=60n nw=240n
XXI9 c cn net46 net099 VDD VSS / TG pl=60n pw=340n nl=60n nw=240n
XXI32 cn c net076 net33 VDD VSS / TG pl=60n pw=260n nl=60n nw=200n
XXI34 SE VDD VSS SEN / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net099 VDD VSS QN / INV pl=60n pw=400n nl=60n nw=280n
XXI31 RN VDD VSS r / INV pl=60n pw=280n nl=60n nw=200n
XXI5 net0147 VDD VSS Q / INV pl=60n pw=400n nl=60n nw=280n
XXI13 c VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net099 VDD VSS net0147 / INV pl=60n pw=320n nl=60n nw=260n
XXI4 CKN VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFNRX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFNRX3H7L CKN D Q QN RN SE SI VDD VSS
*.PININFO CKN:I D:I RN:I SE:I SI:I Q:O QN:O VDD:B VSS:B
XXI32 cn c net076 net33 VDD VSS / TG pl=60n pw=360n nl=60n nw=260n
XXI9 c cn net46 net099 VDD VSS / TG pl=60n pw=360n nl=60n nw=260n
XXI4 CKN VDD VSS c / INV pl=60n pw=340n nl=60n nw=240n
XXI10 net099 VDD VSS net0147 / INV pl=60n pw=360n nl=60n nw=260n
XXI13 c VDD VSS cn / INV pl=60n pw=340n nl=60n nw=240n
XXI5 net0147 VDD VSS Q / INV pl=60n pw=600n nl=60n nw=420n
XXI31 RN VDD VSS r / INV pl=60n pw=340n nl=60n nw=240n
XXI12 net099 VDD VSS QN / INV pl=60n pw=600n nl=60n nw=420n
XXI34 SE VDD VSS SEN / INV pl=60n pw=340n nl=60n nw=240n
MMN1 net099 cn net53 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net53 net0147 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net099 r VSS VSS nm1p2_lvt_lp W=260n L=60n m=1
MMN4 net46 net33 VSS VSS nm1p2_lvt_lp W=260n L=60n m=1
MMP4 net54 r VDD VDD pm1p2_lvt_lp W=360n L=60n m=1
MMP2 net48 net0147 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net099 c net48 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=360n L=60n m=1
XXI30 D SEN SE VDD VSS net076 / TSINV pl=60n pw=340n nl=60n nw=260n
XXI33 SI SE SEN VDD VSS net076 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI29 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFNSRX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFNSRX0P5H7L CKN D Q QN RN SE SI SN VDD VSS
*.PININFO CKN:I D:I RN:I SE:I SI:I SN:I Q:O QN:O VDD:B VSS:B
MMN5 net062 SN VSS VSS nm1p2_lvt_lp W=220n L=60n m=1
MMN1 net0115 cn net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0167 net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN6 net0115 r net062 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN4 net46 net33 net062 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMP4 net0115 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP5 net54 r VDD VDD pm1p2_lvt_lp W=280n L=60n m=1
MMP2 net67 net0167 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net0115 c net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=300n L=60n m=1
XXI29 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI33 SI SE SEN VDD VSS net087 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI30 D SEN SE VDD VSS net087 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI35 cn c net087 net33 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
XXI9 c cn net46 net0115 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
XI3 RN VDD VSS r / INV pl=60n pw=280n nl=60n nw=200n
XI1 c VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
XI2 SE VDD VSS SEN / INV pl=60n pw=280n nl=60n nw=200n
XI0 CKN VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net0115 VDD VSS QN / INV pl=60n pw=280n nl=60n nw=200n
XXI5 net0167 VDD VSS Q / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net0115 VDD VSS net0167 / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFNSRX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFNSRX1H7L CKN D Q QN RN SE SI SN VDD VSS
*.PININFO CKN:I D:I RN:I SE:I SI:I SN:I Q:O QN:O VDD:B VSS:B
MNM4 net46 net33 net062 VSS nm1p2_lvt_lp W=220n L=60n m=1
MNM3 net0115 r net062 VSS nm1p2_lvt_lp W=200n L=60n m=1
MNM2 net76 net0167 net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net0115 cn net76 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net062 SN VSS VSS nm1p2_lvt_lp W=220n L=60n m=1
MPM4 net46 net33 net54 VDD pm1p2_lvt_lp W=300n L=60n m=1
MPM3 net0115 c net79 VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM2 net79 net0167 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM1 net54 r VDD VDD pm1p2_lvt_lp W=300n L=60n m=1
MPM0 net0115 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
XI0 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI33 SI SE SEN VDD VSS net087 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI30 D SEN SE VDD VSS net087 / TSINV pl=60n pw=280n nl=60n nw=200n
XI4 c cn net46 net0115 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
XXI35 cn c net087 net33 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
XI8 CKN VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XI7 c VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
XI6 SE VDD VSS SEN / INV pl=60n pw=280n nl=60n nw=200n
XI5 RN VDD VSS r / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net0115 VDD VSS QN / INV pl=60n pw=340n nl=60n nw=240n
XXI5 net0167 VDD VSS Q / INV pl=60n pw=340n nl=60n nw=240n
XXI10 net0115 VDD VSS net0167 / INV pl=60n pw=300n nl=60n nw=220n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFNSX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFNSX0P5H7L CKN D Q QN SE SI SN VDD VSS
*.PININFO CKN:I D:I SE:I SI:I SN:I Q:O QN:O VDD:B VSS:B
MMN6 net056 SN VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN1 net0100 cn net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net048 net056 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 net056 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMP0 net0100 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP2 net67 net048 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net0100 c net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 VDD VDD pm1p2_lvt_lp W=280n L=60n m=1
XXI32 SI SE SEN VDD VSS net076 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI29 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI30 D SEN SE VDD VSS net076 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI9 c cn net46 net0100 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
XXI33 cn c net076 net33 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
XXI34 SE VDD VSS SEN / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net0100 VDD VSS QN / INV pl=60n pw=280n nl=60n nw=200n
XXI5 net048 VDD VSS Q / INV pl=60n pw=280n nl=60n nw=200n
XXI13 c VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net0100 VDD VSS net048 / INV pl=60n pw=280n nl=60n nw=200n
XXI4 CKN VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFNSX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFNSX1H7L CKN D Q QN SE SI SN VDD VSS
*.PININFO CKN:I D:I SE:I SI:I SN:I Q:O QN:O VDD:B VSS:B
MMN6 net056 SN VSS VSS nm1p2_lvt_lp W=220n L=60n m=1
MMN1 net0100 cn net26 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net26 net048 net056 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 net056 VSS nm1p2_lvt_lp W=220n L=60n m=1
MMP0 net0100 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP2 net67 net048 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net0100 c net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 VDD VDD pm1p2_lvt_lp W=300n L=60n m=1
XXI32 SI SE SEN VDD VSS net076 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI29 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI30 D SEN SE VDD VSS net076 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI9 c cn net46 net0100 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
XXI33 cn c net076 net33 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
XXI34 SE VDD VSS SEN / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net0100 VDD VSS QN / INV pl=60n pw=340n nl=60n nw=240n
XXI5 net048 VDD VSS Q / INV pl=60n pw=340n nl=60n nw=240n
XXI13 c VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net0100 VDD VSS net048 / INV pl=60n pw=300n nl=60n nw=220n
XXI4 CKN VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFNSX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFNSX2H7L CKN D Q QN SE SI SN VDD VSS
*.PININFO CKN:I D:I SE:I SI:I SN:I Q:O QN:O VDD:B VSS:B
MMN6 net056 SN VSS VSS nm1p2_lvt_lp W=240n L=60n m=1
MMN1 net0100 cn net26 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net26 net048 net056 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 net056 VSS nm1p2_lvt_lp W=240n L=60n m=1
MMP0 net0100 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP2 net67 net048 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net0100 c net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 VDD VDD pm1p2_lvt_lp W=340n L=60n m=1
XXI32 SI SE SEN VDD VSS net076 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI29 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI30 D SEN SE VDD VSS net076 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI9 c cn net46 net0100 VDD VSS / TG pl=60n pw=340n nl=60n nw=240n
XXI33 cn c net076 net33 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
XXI34 SE VDD VSS SEN / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net0100 VDD VSS QN / INV pl=60n pw=400n nl=60n nw=280n
XXI5 net048 VDD VSS Q / INV pl=60n pw=400n nl=60n nw=280n
XXI13 c VDD VSS cn / INV pl=60n pw=340n nl=60n nw=240n
XXI10 net0100 VDD VSS net048 / INV pl=60n pw=340n nl=60n nw=240n
XXI4 CKN VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFNX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFNX0P5H7L CKN D Q QN SE SI VDD VSS
*.PININFO CKN:I D:I SE:I SI:I Q:O QN:O VDD:B VSS:B
XXI9 net44 net42 net69 VDD VSS net51 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI21 D net56 SE VDD VSS net76 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI22 SI SE net56 VDD VSS net76 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI15 net48 net69 net42 VDD VSS net51 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI14 net44 net42 net69 VDD VSS net39 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI23 SE VDD VSS net56 / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net51 VDD VSS net48 / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net51 VDD VSS Q / INV pl=60n pw=280n nl=60n nw=200n
XXI4 CKN VDD VSS net42 / INV pl=60n pw=280n nl=60n nw=200n
XXI5 net48 VDD VSS QN / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net39 VDD VSS net44 / INV pl=60n pw=280n nl=60n nw=200n
XXI13 net42 VDD VSS net69 / INV pl=60n pw=280n nl=60n nw=200n
XXI6 net69 net42 net76 net39 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFNX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFNX1H7L CKN D Q QN SE SI VDD VSS
*.PININFO CKN:I D:I SE:I SI:I Q:O QN:O VDD:B VSS:B
XXI9 net44 net42 net69 VDD VSS net51 / TSINV pl=60n pw=300n nl=60n nw=220n
XXI21 D net56 SE VDD VSS net76 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI22 SI SE net56 VDD VSS net76 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI15 net48 net69 net42 VDD VSS net51 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI14 net44 net42 net69 VDD VSS net39 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI23 SE VDD VSS net56 / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net51 VDD VSS net48 / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net51 VDD VSS Q / INV pl=60n pw=340n nl=60n nw=240n
XXI4 CKN VDD VSS net42 / INV pl=60n pw=280n nl=60n nw=200n
XXI5 net48 VDD VSS QN / INV pl=60n pw=340n nl=60n nw=240n
XXI7 net39 VDD VSS net44 / INV pl=60n pw=300n nl=60n nw=220n
XXI13 net42 VDD VSS net69 / INV pl=60n pw=280n nl=60n nw=200n
XXI6 net69 net42 net76 net39 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFNX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFNX2H7L CKN D Q QN SE SI VDD VSS
*.PININFO CKN:I D:I SE:I SI:I Q:O QN:O VDD:B VSS:B
XXI21 D net56 SE VDD VSS net76 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI22 SI SE net56 VDD VSS net76 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI15 net48 net69 net42 VDD VSS net51 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI14 net44 net42 net69 VDD VSS net39 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI9 net44 net42 net69 VDD VSS net51 / TSINV pl=60n pw=340n nl=60n nw=240n
XXI23 SE VDD VSS net56 / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net51 VDD VSS Q / INV pl=60n pw=400n nl=60n nw=280n
XXI10 net51 VDD VSS net48 / INV pl=60n pw=280n nl=60n nw=200n
XXI4 CKN VDD VSS net42 / INV pl=60n pw=280n nl=60n nw=200n
XXI13 net42 VDD VSS net69 / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net39 VDD VSS net44 / INV pl=60n pw=340n nl=60n nw=240n
XXI5 net48 VDD VSS QN / INV pl=60n pw=400n nl=60n nw=280n
XXI6 net69 net42 net76 net39 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFNX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFNX3H7L CKN D Q QN SE SI VDD VSS
*.PININFO CKN:I D:I SE:I SI:I Q:O QN:O VDD:B VSS:B
XXI6 net69 net42 net76 net39 VDD VSS / TG pl=60n pw=340n nl=60n nw=240n
XXI5 net48 VDD VSS QN / INV pl=60n pw=600n nl=60n nw=420n
XXI7 net39 VDD VSS net44 / INV pl=60n pw=360n nl=60n nw=260n
XXI13 net42 VDD VSS net69 / INV pl=60n pw=340n nl=60n nw=240n
XXI4 CKN VDD VSS net42 / INV pl=60n pw=340n nl=60n nw=240n
XXI10 net51 VDD VSS net48 / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net51 VDD VSS Q / INV pl=60n pw=600n nl=60n nw=420n
XXI23 SE VDD VSS net56 / INV pl=60n pw=340n nl=60n nw=240n
XXI22 SI SE net56 VDD VSS net76 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI15 net48 net69 net42 VDD VSS net51 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI14 net44 net42 net69 VDD VSS net39 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI9 net44 net42 net69 VDD VSS net51 / TSINV pl=60n pw=360n nl=60n nw=260n
XXI21 D net56 SE VDD VSS net76 / TSINV pl=60n pw=340n nl=60n nw=240n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFQX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFQX0P5H7L CK D Q SE SI VDD VSS
*.PININFO CK:I D:I SE:I SI:I Q:O VDD:B VSS:B
XXI14 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI18 SI SE sen VDD VSS net050 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI16 D sen SE VDD VSS net050 / TSINV pl=60n pw=300n nl=60n nw=220n
XXI9 net46 c cn VDD VSS net25 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI15 net9 cn c VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI19 SE VDD VSS sen / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=280n nl=60n nw=200n
XXI13 cn VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net25 VDD VSS Q / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XXI4 CK VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
XXI17 cn c net050 net33 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFQX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFQX1H7L CK D Q SE SI VDD VSS
*.PININFO CK:I D:I SE:I SI:I Q:O VDD:B VSS:B
XXI15 net9 cn c VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI9 net46 c cn VDD VSS net25 / TSINV pl=60n pw=300n nl=60n nw=220n
XXI16 D sen SE VDD VSS net050 / TSINV pl=60n pw=300n nl=60n nw=220n
XXI18 SI SE sen VDD VSS net050 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI14 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI4 CK VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net25 VDD VSS Q / INV pl=60n pw=340n nl=60n nw=240n
XXI13 cn VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=300n nl=60n nw=220n
XXI19 SE VDD VSS sen / INV pl=60n pw=280n nl=60n nw=200n
XXI17 cn c net050 net33 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFQX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFQX2H7L CK D Q SE SI VDD VSS
*.PININFO CK:I D:I SE:I SI:I Q:O VDD:B VSS:B
XXI16 D sen SE VDD VSS net050 / TSINV pl=60n pw=300n nl=60n nw=220n
XXI15 net9 cn c VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI9 net46 c cn VDD VSS net25 / TSINV pl=60n pw=340n nl=60n nw=240n
XXI18 SI SE sen VDD VSS net050 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI14 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI13 cn VDD VSS c / INV pl=60n pw=340n nl=60n nw=240n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=340n nl=60n nw=240n
XXI19 SE VDD VSS sen / INV pl=60n pw=340n nl=60n nw=240n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net25 VDD VSS Q / INV pl=60n pw=400n nl=60n nw=280n
XXI4 CK VDD VSS cn / INV pl=60n pw=340n nl=60n nw=240n
XXI17 cn c net050 net33 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFQX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFQX3H7L CK D Q SE SI VDD VSS
*.PININFO CK:I D:I SE:I SI:I Q:O VDD:B VSS:B
XXI4 CK VDD VSS cn / INV pl=60n pw=340n nl=60n nw=240n
XXI12 net25 VDD VSS Q / INV pl=60n pw=600n nl=60n nw=420n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XXI19 SE VDD VSS sen / INV pl=60n pw=340n nl=60n nw=240n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=360n nl=60n nw=260n
XXI13 cn VDD VSS c / INV pl=60n pw=340n nl=60n nw=240n
XXI17 cn c net050 net33 VDD VSS / TG pl=60n pw=340n nl=60n nw=240n
XXI14 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI18 SI SE sen VDD VSS net050 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI9 net46 c cn VDD VSS net25 / TSINV pl=60n pw=360n nl=60n nw=260n
XXI15 net9 cn c VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI16 D sen SE VDD VSS net050 / TSINV pl=60n pw=340n nl=60n nw=240n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFRQX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFRQX0P5H7L CK D Q RN SE SI VDD VSS
*.PININFO CK:I D:I RN:I SE:I SI:I Q:O VDD:B VSS:B
XXI9 c cn net46 net0182 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
XXI12 net0182 VDD VSS Q / INV pl=60n pw=280n nl=60n nw=200n
XXI32 SE VDD VSS sen / INV pl=60n pw=280n nl=60n nw=200n
XXI4 CK VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net0182 VDD VSS net048 / INV pl=60n pw=280n nl=60n nw=240n
XXI13 cn VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XXI33 D sen SE VDD VSS net075 / TSINV pl=60n pw=280n nl=60n nw=240n
XXI30 net075 cn c VDD VSS net33 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI29 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI34 SI SE sen VDD VSS net075 / TSINV pl=60n pw=250n nl=60n nw=200n
MMP1 net0182 c net062 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP2 net062 net048 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP0 net0182 RN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP3 net46 net33 VDD VDD pm1p2_lvt_lp W=280n L=60n m=1
MMN1 net0182 cn net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN6 net056 RN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 net056 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN2 net36 net048 net056 VSS nm1p2_lvt_lp W=150n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFRQX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFRQX1H7L CK D Q RN SE SI VDD VSS
*.PININFO CK:I D:I RN:I SE:I SI:I Q:O VDD:B VSS:B
MMN6 net056 RN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 net0182 cn net25 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net25 net048 net056 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 net056 VSS nm1p2_lvt_lp W=220n L=60n m=1
MMP0 net0182 RN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP2 net062 net048 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net0182 c net062 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 VDD VDD pm1p2_lvt_lp W=300n L=60n m=1
XXI33 D sen SE VDD VSS net075 / TSINV pl=60n pw=280n nl=60n nw=240n
XXI34 SI SE sen VDD VSS net075 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI29 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI30 net075 cn c VDD VSS net33 / TSINV pl=60n pw=300n nl=60n nw=220n
XXI32 SE VDD VSS sen / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net0182 VDD VSS Q / INV pl=60n pw=340n nl=60n nw=240n
XXI13 cn VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net0182 VDD VSS net048 / INV pl=60n pw=280n nl=60n nw=240n
XXI4 CK VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
XXI9 c cn net46 net0182 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFRQX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFRQX2H7L CK D Q RN SE SI VDD VSS
*.PININFO CK:I D:I RN:I SE:I SI:I Q:O VDD:B VSS:B
MMN6 net056 RN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 net0182 cn net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net048 net056 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 net056 VSS nm1p2_lvt_lp W=240n L=60n m=1
MMP0 net0182 RN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP2 net062 net048 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net0182 c net062 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 VDD VDD pm1p2_lvt_lp W=340n L=60n m=1
XXI33 D sen SE VDD VSS net075 / TSINV pl=60n pw=280n nl=60n nw=240n
XXI34 SI SE sen VDD VSS net075 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI29 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI30 net075 cn c VDD VSS net33 / TSINV pl=60n pw=340n nl=60n nw=240n
XXI32 SE VDD VSS sen / INV pl=60n pw=340n nl=60n nw=240n
XXI12 net0182 VDD VSS Q / INV pl=60n pw=400n nl=60n nw=280n
XXI13 cn VDD VSS c / INV pl=60n pw=340n nl=60n nw=240n
XXI10 net0182 VDD VSS net048 / INV pl=60n pw=280n nl=60n nw=240n
XXI4 CK VDD VSS cn / INV pl=60n pw=340n nl=60n nw=240n
XXI9 c cn net46 net0182 VDD VSS / TG pl=60n pw=340n nl=60n nw=240n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFRQX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFRQX3H7L CK D Q RN SE SI VDD VSS
*.PININFO CK:I D:I RN:I SE:I SI:I Q:O VDD:B VSS:B
MNM3 net056 RN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM2 net0182 cn net89 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net89 net048 net056 VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net46 net33 net056 VSS nm1p2_lvt_lp W=260n L=60n m=1
MPM0 net46 net33 VDD VDD pm1p2_lvt_lp W=360n L=60n m=1
MPM3 net0182 RN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MPM2 net84 net048 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM1 net0182 c net84 VDD pm1p2_lvt_lp W=150n L=60n m=1
XI3 D sen SE VDD VSS net075 / TSINV pl=60n pw=320n nl=60n nw=240n
XI2 SI SE sen VDD VSS net075 / TSINV pl=60n pw=250n nl=60n nw=200n
XI1 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XI0 net075 cn c VDD VSS net33 / TSINV pl=60n pw=360n nl=60n nw=260n
XXI12 net0182 VDD VSS Q / INV pl=60n pw=600n nl=60n nw=420n
XXI10 net0182 VDD VSS net048 / INV pl=60n pw=600n nl=60n nw=420n
XI8 SE VDD VSS sen / INV pl=60n pw=340n nl=60n nw=240n
XI4 CK VDD VSS cn / INV pl=60n pw=340n nl=60n nw=240n
XI6 cn VDD VSS c / INV pl=60n pw=340n nl=60n nw=240n
XI9 c cn net46 net0182 VDD VSS / TG pl=60n pw=360n nl=60n nw=260n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFRX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFRX0P5H7L CK D Q QN RN SE SI VDD VSS
*.PININFO CK:I D:I RN:I SE:I SI:I Q:O QN:O VDD:B VSS:B
MMN1 net099 cn net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0146 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net099 r VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMP4 net54 r VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP2 net67 net0146 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net099 c net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=280n L=60n m=1
XXI29 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI33 SI SE sen VDD VSS net076 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI30 D sen SE VDD VSS net076 / TSINV pl=60n pw=280n nl=60n nw=240n
XXI9 c cn net46 net099 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
XXI32 cn c net076 net33 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
XXI34 SE VDD VSS sen / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net099 VDD VSS QN / INV pl=60n pw=280n nl=60n nw=200n
XXI31 RN VDD VSS r / INV pl=60n pw=280n nl=60n nw=200n
XXI5 net0146 VDD VSS Q / INV pl=60n pw=280n nl=60n nw=200n
XXI13 cn VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net099 VDD VSS net0146 / INV pl=60n pw=280n nl=60n nw=240n
XXI4 CK VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFRX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFRX1H7L CK D Q QN RN SE SI VDD VSS
*.PININFO CK:I D:I RN:I SE:I SI:I Q:O QN:O VDD:B VSS:B
MNM3 net46 net33 VSS VSS nm1p2_lvt_lp W=220n L=60n m=1
MNM2 net099 r VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 net35 net0146 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM0 net099 cn net35 VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM3 net46 net33 net54 VDD pm1p2_lvt_lp W=300n L=60n m=1
MPM2 net099 c net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM1 net67 net0146 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MPM0 net54 r VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
XI2 D sen SE VDD VSS net076 / TSINV pl=60n pw=280n nl=60n nw=240n
XI1 SI SE sen VDD VSS net076 / TSINV pl=60n pw=250n nl=60n nw=200n
XI0 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XI4 cn c net076 net33 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
XI3 c cn net46 net099 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
XI11 CK VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
XI10 net099 VDD VSS net0146 / INV pl=60n pw=280n nl=60n nw=240n
XI9 cn VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XI8 net0146 VDD VSS Q / INV pl=60n pw=340n nl=60n nw=240n
XI7 RN VDD VSS r / INV pl=60n pw=280n nl=60n nw=200n
XI6 net099 VDD VSS QN / INV pl=60n pw=340n nl=60n nw=240n
XI5 SE VDD VSS sen / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net15 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 net15 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP2 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFRX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFRX2H7L CK D Q QN RN SE SI VDD VSS
*.PININFO CK:I D:I RN:I SE:I SI:I Q:O QN:O VDD:B VSS:B
MMN0 net55 cn net43 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net40 RN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 net43 net41 net40 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP2 net55 RN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP0 net55 c net059 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net059 net41 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
XXI29 SI SE sen VDD VSS net77 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI28 D sen SE VDD VSS net77 / TSINV pl=60n pw=280n nl=60n nw=240n
XXI21 net66 c cn VDD VSS net61 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI6 net77 cn c VDD VSS net61 / TSINV pl=60n pw=340n nl=60n nw=240n
XXI32 net61 RN VDD VSS net66 / NAND2 pl=60n pw=340n nl=60n nw=240n
XXI27 net41 VDD VSS QN / INV pl=60n pw=400n nl=60n nw=280n
XXI19 net55 VDD VSS net41 / INV pl=60n pw=280n nl=60n nw=240n
XXI13 cn VDD VSS c / INV pl=60n pw=340n nl=60n nw=240n
XXI30 SE VDD VSS sen / INV pl=60n pw=340n nl=60n nw=240n
XXI26 net55 VDD VSS Q / INV pl=60n pw=400n nl=60n nw=280n
XXI4 CK VDD VSS cn / INV pl=60n pw=340n nl=60n nw=240n
XXI22 c cn net66 net55 VDD VSS / TG pl=60n pw=340n nl=60n nw=240n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net15 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 net15 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP2 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFRX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFRX3H7L CK D Q QN RN SE SI VDD VSS
*.PININFO CK:I D:I RN:I SE:I SI:I Q:O QN:O VDD:B VSS:B
XXI4 CK VDD VSS cn / INV pl=60n pw=340n nl=60n nw=240n
XXI26 net55 VDD VSS Q / INV pl=60n pw=600n nl=60n nw=420n
XXI30 SE VDD VSS sen / INV pl=60n pw=340n nl=60n nw=240n
XXI13 cn VDD VSS c / INV pl=60n pw=340n nl=60n nw=240n
XXI19 net55 VDD VSS net41 / INV pl=60n pw=360n nl=60n nw=260n
XXI27 net41 VDD VSS QN / INV pl=60n pw=600n nl=60n nw=420n
XXI22 c cn net66 net55 VDD VSS / TG pl=60n pw=360n nl=60n nw=260n
MMN0 net55 cn net43 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net17 RN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 net43 net41 net17 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMP2 net55 RN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP0 net55 c net26 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net26 net41 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
XXI32 net61 RN VDD VSS net66 / NAND2 pl=60n pw=360n nl=60n nw=260n
XXI6 net77 cn c VDD VSS net61 / TSINV pl=60n pw=360n nl=60n nw=260n
XXI21 net66 c cn VDD VSS net61 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI28 D sen SE VDD VSS net77 / TSINV pl=60n pw=320n nl=60n nw=240n
XXI29 SI SE sen VDD VSS net77 / TSINV pl=60n pw=250n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFSQX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFSQX1H7L CK D Q SE SI SN VDD VSS
*.PININFO CK:I D:I SE:I SI:I SN:I Q:O VDD:B VSS:B
MMN1 net0187 cn net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net048 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net0187 s VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net087 net33 VSS VSS nm1p2_lvt_lp W=190n L=60n m=1
MMP4 net54 s VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP2 net068 net048 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net0187 c net068 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net087 net33 net54 VDD pm1p2_lvt_lp W=170n L=60n m=1
XXI35 SI SE sen VDD VSS net080 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI34 D sen SE VDD VSS net080 / TSINV pl=60n pw=250n nl=60n nw=180n
XXI29 net087 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI30 net080 cn c VDD VSS net33 / TSINV pl=60n pw=190n nl=60n nw=190n
XXI33 SE VDD VSS sen / INV pl=60n pw=210n nl=60n nw=170n
XXI12 net0187 VDD VSS Q / INV pl=60n pw=270n nl=60n nw=210n
XXI31 SN VDD VSS s / INV pl=60n pw=210n nl=60n nw=170n
XXI13 cn VDD VSS c / INV pl=60n pw=210n nl=60n nw=170n
XXI10 net0187 VDD VSS net048 / INV pl=60n pw=190n nl=60n nw=150n
XXI4 CK VDD VSS cn / INV pl=60n pw=210n nl=60n nw=170n
XXI9 c cn net087 net0187 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFSQX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFSQX2H7L CK D Q SE SI SN VDD VSS
*.PININFO CK:I D:I SE:I SI:I SN:I Q:O VDD:B VSS:B
MMN1 net0187 cn net29 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net29 net048 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net0187 s VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net087 net33 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMP4 net54 s VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP2 net068 net048 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net0187 c net068 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net087 net33 net54 VDD pm1p2_lvt_lp W=180n L=60n m=1
XXI35 SI SE sen VDD VSS net080 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI34 D sen SE VDD VSS net080 / TSINV pl=60n pw=270n nl=60n nw=190n
XXI29 net087 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI30 net080 cn c VDD VSS net33 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI33 SE VDD VSS sen / INV pl=60n pw=210n nl=60n nw=170n
XXI12 net0187 VDD VSS Q / INV pl=60n pw=380n nl=60n nw=300n
XXI31 SN VDD VSS s / INV pl=60n pw=210n nl=60n nw=170n
XXI13 cn VDD VSS c / INV pl=60n pw=210n nl=60n nw=170n
XXI10 net0187 VDD VSS net048 / INV pl=60n pw=190n nl=60n nw=150n
XXI4 CK VDD VSS cn / INV pl=60n pw=210n nl=60n nw=170n
XXI9 c cn net087 net0187 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFSQX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFSQX3H7L CK D Q SE SI SN VDD VSS
*.PININFO CK:I D:I SE:I SI:I SN:I Q:O VDD:B VSS:B
MMP3 net087 net33 net54 VDD pm1p2_lvt_lp W=180n L=60n m=1
MMP1 net0187 c net068 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP4 net54 s VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP2 net068 net048 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
XXI33 SE VDD VSS sen / INV pl=60n pw=210n nl=60n nw=170n
XXI4 CK VDD VSS cn / INV pl=60n pw=210n nl=60n nw=170n
XXI10 net0187 VDD VSS net048 / INV pl=60n pw=250n nl=60n nw=200n
XXI12 net0187 VDD VSS Q / INV pl=60n pw=570n nl=60n nw=450n
XXI31 SN VDD VSS s / INV pl=60n pw=210n nl=60n nw=170n
XXI13 cn VDD VSS c / INV pl=60n pw=210n nl=60n nw=170n
XXI9 c cn net087 net0187 VDD VSS / TG pl=60n pw=250n nl=60n nw=200n
MMN1 net0187 cn net29 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net29 net048 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net0187 s VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net087 net33 VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
XXI35 SI SE sen VDD VSS net080 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI30 net080 cn c VDD VSS net33 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI29 net087 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI34 D sen SE VDD VSS net080 / TSINV pl=60n pw=270n nl=60n nw=190n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFSRQX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFSRQX1H7L CK D Q RN SE SI SN VDD VSS
*.PININFO CK:I D:I RN:I SE:I SI:I SN:I Q:O VDD:B VSS:B
MMN5 net062 SN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 net0115 cn net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net093 net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN6 net0115 r net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 net062 VSS nm1p2_lvt_lp W=190n L=60n m=1
MMP4 net0115 SN VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP5 net54 r VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP2 net67 net093 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net0115 c net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=170n L=60n m=1
XXI33 SI SE sen VDD VSS net088 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI29 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI30 D sen SE VDD VSS net088 / TSINV pl=60n pw=250n nl=60n nw=180n
XXI35 cn c net088 net33 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI9 c cn net46 net0115 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI32 RN VDD VSS r / INV pl=60n pw=210n nl=60n nw=170n
XXI34 SE VDD VSS sen / INV pl=60n pw=210n nl=60n nw=170n
XXI5 net093 VDD VSS Q / INV pl=60n pw=270n nl=60n nw=210n
XXI13 cn VDD VSS c / INV pl=60n pw=210n nl=60n nw=170n
XXI10 net0115 VDD VSS net093 / INV pl=60n pw=190n nl=60n nw=150n
XXI4 CK VDD VSS cn / INV pl=60n pw=210n nl=60n nw=170n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFSRQX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFSRQX2H7L CK D Q RN SE SI SN VDD VSS
*.PININFO CK:I D:I RN:I SE:I SI:I SN:I Q:O VDD:B VSS:B
MMN5 net062 SN VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 net0115 cn net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net093 net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN6 net0115 r net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 net062 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMP4 net0115 SN VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP5 net54 r VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP2 net67 net093 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net0115 c net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=180n L=60n m=1
XXI33 SI SE sen VDD VSS net088 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI29 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI30 D sen SE VDD VSS net088 / TSINV pl=60n pw=270n nl=60n nw=190n
XXI35 cn c net088 net33 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI9 c cn net46 net0115 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI32 RN VDD VSS r / INV pl=60n pw=210n nl=60n nw=170n
XXI34 SE VDD VSS sen / INV pl=60n pw=210n nl=60n nw=170n
XXI5 net093 VDD VSS Q / INV pl=60n pw=380n nl=60n nw=300n
XXI13 cn VDD VSS c / INV pl=60n pw=210n nl=60n nw=170n
XXI10 net0115 VDD VSS net093 / INV pl=60n pw=210n nl=60n nw=170n
XXI4 CK VDD VSS cn / INV pl=60n pw=210n nl=60n nw=170n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFSRQX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFSRQX3H7L CK D Q RN SE SI SN VDD VSS
*.PININFO CK:I D:I RN:I SE:I SI:I SN:I Q:O VDD:B VSS:B
XXI9 c cn net46 net0115 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI35 cn c net088 net33 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI4 CK VDD VSS cn / INV pl=60n pw=210n nl=60n nw=170n
XXI10 net0115 VDD VSS net093 / INV pl=60n pw=250n nl=60n nw=200n
XXI13 cn VDD VSS c / INV pl=60n pw=210n nl=60n nw=170n
XXI5 net093 VDD VSS Q / INV pl=60n pw=570n nl=60n nw=450n
XXI34 SE VDD VSS sen / INV pl=60n pw=210n nl=60n nw=170n
XXI32 RN VDD VSS r / INV pl=60n pw=210n nl=60n nw=170n
MMN5 net062 SN VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN1 net0115 cn net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net093 net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN6 net0115 r net062 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN4 net46 net33 net062 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMP4 net0115 SN VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP5 net54 r VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP2 net67 net093 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net0115 c net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=180n L=60n m=1
XXI30 D sen SE VDD VSS net088 / TSINV pl=60n pw=270n nl=60n nw=190n
XXI29 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI33 SI SE sen VDD VSS net088 / TSINV pl=60n pw=150n nl=60n nw=150n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFSRX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFSRX0P5H7L CK D Q QN RN SE SI SN VDD VSS
*.PININFO CK:I D:I RN:I SE:I SI:I SN:I Q:O QN:O VDD:B VSS:B
MMN5 net062 SN VSS VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN1 net0115 cn net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0164 net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN6 net0115 r net062 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN4 net46 net33 net062 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMP4 net0115 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP5 net54 r VDD VDD pm1p2_lvt_lp W=280n L=60n m=1
MMP2 net67 net0164 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net0115 c net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=280n L=60n m=1
XXI29 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI33 SI SE SEN VDD VSS net087 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI30 D SEN SE VDD VSS net087 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI35 cn c net087 net33 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
XXI9 c cn net46 net0115 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
XXI12 net0115 VDD VSS QN / INV pl=60n pw=280n nl=60n nw=200n
XXI32 RN VDD VSS r / INV pl=60n pw=280n nl=60n nw=200n
XXI34 SE VDD VSS SEN / INV pl=60n pw=280n nl=60n nw=200n
XXI5 net0164 VDD VSS Q / INV pl=60n pw=280n nl=60n nw=200n
XXI13 cn VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net0115 VDD VSS net0164 / INV pl=60n pw=280n nl=60n nw=200n
XXI4 CK VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFSRX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFSRX1H7L CK D Q QN RN SE SI SN VDD VSS
*.PININFO CK:I D:I RN:I SE:I SI:I SN:I Q:O QN:O VDD:B VSS:B
MMN5 net062 SN VSS VSS nm1p2_lvt_lp W=220n L=60n m=1
MMN1 net0115 cn net35 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net35 net0164 net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN6 net0115 r net062 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN4 net46 net33 net062 VSS nm1p2_lvt_lp W=220n L=60n m=1
MMP4 net0115 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP5 net54 r VDD VDD pm1p2_lvt_lp W=300n L=60n m=1
MMP2 net67 net0164 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net0115 c net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=300n L=60n m=1
XXI29 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI33 SI SE SEN VDD VSS net087 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI30 D SEN SE VDD VSS net087 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI35 cn c net087 net33 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
XXI9 c cn net46 net0115 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
XXI12 net0115 VDD VSS QN / INV pl=60n pw=280n nl=60n nw=200n
XXI32 RN VDD VSS r / INV pl=60n pw=280n nl=60n nw=200n
XXI34 SE VDD VSS SEN / INV pl=60n pw=280n nl=60n nw=200n
XXI5 net0164 VDD VSS Q / INV pl=60n pw=280n nl=60n nw=200n
XXI13 cn VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net0115 VDD VSS net0164 / INV pl=60n pw=300n nl=60n nw=220n
XXI4 CK VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFSRX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFSRX2H7L CK D Q QN RN SE SI SN VDD VSS
*.PININFO CK:I D:I RN:I SE:I SI:I SN:I Q:O QN:O VDD:B VSS:B
MMN4 net46 net33 net062 VSS nm1p2_lvt_lp W=240n L=60n m=1
MMN6 net0115 r net062 VSS nm1p2_lvt_lp W=200n L=60n m=1
MMN2 net35 net0164 net062 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN1 net0115 cn net35 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN5 net062 SN VSS VSS nm1p2_lvt_lp W=240n L=60n m=1
MMP3 net46 net33 net54 VDD pm1p2_lvt_lp W=340n L=60n m=1
MMP1 net0115 c net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP2 net67 net0164 net54 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP5 net54 r VDD VDD pm1p2_lvt_lp W=340n L=60n m=1
MMP4 net0115 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
XXI30 D SEN SE VDD VSS net087 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI33 SI SE SEN VDD VSS net087 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI29 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI9 c cn net46 net0115 VDD VSS / TG pl=60n pw=340n nl=60n nw=240n
XXI35 cn c net087 net33 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
XXI4 CK VDD VSS cn / INV pl=60n pw=340n nl=60n nw=240n
XXI10 net0115 VDD VSS net0164 / INV pl=60n pw=340n nl=60n nw=240n
XXI13 cn VDD VSS c / INV pl=60n pw=340n nl=60n nw=240n
XXI5 net0164 VDD VSS Q / INV pl=60n pw=400n nl=60n nw=280n
XXI34 SE VDD VSS SEN / INV pl=60n pw=340n nl=60n nw=240n
XXI32 RN VDD VSS r / INV pl=60n pw=340n nl=60n nw=240n
XXI12 net0115 VDD VSS QN / INV pl=60n pw=400n nl=60n nw=280n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFSX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFSX0P5H7L CK D Q QN SE SI SN VDD VSS
*.PININFO CK:I D:I SE:I SI:I SN:I Q:O QN:O VDD:B VSS:B
MMN6 net056 SN VSS VSS nm1p2_lvt_lp W=240n L=60n m=1
MMN1 net099 cn net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0146 net056 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 net056 VSS nm1p2_lvt_lp W=240n L=60n m=1
MMP0 net099 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP2 net67 net0146 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net099 c net67 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 VDD VDD pm1p2_lvt_lp W=280n L=60n m=1
XXI32 SI SE sen VDD VSS net076 / TSINV pl=60n pw=250n nl=60n nw=180n
XXI29 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI30 D sen SE VDD VSS net076 / TSINV pl=60n pw=280n nl=60n nw=210n
XXI9 c cn net46 net099 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
XXI33 cn c net076 net33 VDD VSS / TG pl=60n pw=300n nl=60n nw=210n
XXI34 SE VDD VSS sen / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net099 VDD VSS QN / INV pl=60n pw=280n nl=60n nw=200n
XXI5 net0146 VDD VSS Q / INV pl=60n pw=280n nl=60n nw=200n
XXI13 cn VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net099 VDD VSS net0146 / INV pl=60n pw=280n nl=60n nw=200n
XXI4 CK VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFSX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFSX1H7L CK D Q QN SE SI SN VDD VSS
*.PININFO CK:I D:I SE:I SI:I SN:I Q:O QN:O VDD:B VSS:B
MMN6 net056 SN VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMN1 net099 cn net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0146 net056 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 net056 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMP0 net099 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP2 net26 net0146 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net099 c net26 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 VDD VDD pm1p2_lvt_lp W=300n L=60n m=1
XXI32 SI SE sen VDD VSS net076 / TSINV pl=60n pw=250n nl=60n nw=180n
XXI29 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI30 D sen SE VDD VSS net076 / TSINV pl=60n pw=280n nl=60n nw=210n
XXI9 c cn net46 net099 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
XXI33 cn c net076 net33 VDD VSS / TG pl=60n pw=300n nl=60n nw=210n
XXI34 SE VDD VSS sen / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net099 VDD VSS QN / INV pl=60n pw=340n nl=60n nw=240n
XXI5 net0146 VDD VSS Q / INV pl=60n pw=340n nl=60n nw=240n
XXI13 cn VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net099 VDD VSS net0146 / INV pl=60n pw=300n nl=60n nw=220n
XXI4 CK VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFSX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFSX2H7L CK D Q QN SE SI SN VDD VSS
*.PININFO CK:I D:I SE:I SI:I SN:I Q:O QN:O VDD:B VSS:B
MMN6 net056 SN VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MMN1 net099 cn net36 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN2 net36 net0146 net056 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN4 net46 net33 net056 VSS nm1p2_lvt_lp W=250n L=60n m=1
MMP0 net099 SN VDD VDD pm1p2_lvt_lp W=200n L=60n m=1
MMP2 net26 net0146 VDD VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP1 net099 c net26 VDD pm1p2_lvt_lp W=150n L=60n m=1
MMP3 net46 net33 VDD VDD pm1p2_lvt_lp W=330n L=60n m=1
XXI32 SI SE sen VDD VSS net076 / TSINV pl=60n pw=250n nl=60n nw=180n
XXI29 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI30 D sen SE VDD VSS net076 / TSINV pl=60n pw=280n nl=60n nw=210n
XXI9 c cn net46 net099 VDD VSS / TG pl=60n pw=340n nl=60n nw=240n
XXI33 cn c net076 net33 VDD VSS / TG pl=60n pw=280n nl=60n nw=210n
XXI34 SE VDD VSS sen / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net099 VDD VSS QN / INV pl=60n pw=400n nl=60n nw=280n
XXI5 net0146 VDD VSS Q / INV pl=60n pw=400n nl=60n nw=280n
XXI13 cn VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net099 VDD VSS net0146 / INV pl=60n pw=340n nl=60n nw=240n
XXI4 CK VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net15 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 net15 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP2 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFTRQX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFTRQX0P5H7L CK D Q RN SE SI VDD VSS
*.PININFO CK:I D:I RN:I SE:I SI:I Q:O VDD:B VSS:B
XXI20 sen SE net034 net046 VDD VSS / TG pl=60n pw=280n nl=60n nw=240n
XXI21 c cn net46 net25 VDD VSS / TG pl=60n pw=280n nl=60n nw=200n
XXI17 D RN VDD VSS net034 / NAND2 pl=60n pw=280n nl=60n nw=240n
XXI15 net9 cn c VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI19 net046 cn c VDD VSS net33 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI22 SI SE sen VDD VSS net046 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI14 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI4 CK VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net25 VDD VSS Q / INV pl=60n pw=280n nl=60n nw=200n
XXI13 cn VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=280n nl=60n nw=200n
XXI23 SE VDD VSS sen / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net15 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 net15 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP2 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFTRQX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFTRQX1H7L CK D Q RN SE SI VDD VSS
*.PININFO CK:I D:I RN:I SE:I SI:I Q:O VDD:B VSS:B
XXI21 c cn net46 net25 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
XXI20 sen SE net034 net046 VDD VSS / TG pl=60n pw=280n nl=60n nw=240n
XXI17 D RN VDD VSS net034 / NAND2 pl=60n pw=280n nl=60n nw=240n
XXI14 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI22 SI SE sen VDD VSS net046 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI19 net046 cn c VDD VSS net33 / TSINV pl=60n pw=300n nl=60n nw=220n
XXI15 net9 cn c VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI23 SE VDD VSS sen / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=300n nl=60n nw=220n
XXI13 cn VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net25 VDD VSS Q / INV pl=60n pw=340n nl=60n nw=240n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=300n nl=60n nw=220n
XXI4 CK VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net15 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 net15 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP2 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFTRQX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFTRQX2H7L CK D Q RN SE SI VDD VSS
*.PININFO CK:I D:I RN:I SE:I SI:I Q:O VDD:B VSS:B
XI1 sen SE net034 net046 VDD VSS / TG pl=60n pw=280n nl=60n nw=240n
XI0 c cn net46 net25 VDD VSS / TG pl=60n pw=340n nl=60n nw=240n
XI2 D RN VDD VSS net034 / NAND2 pl=60n pw=280n nl=60n nw=240n
XI6 net9 cn c VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XI5 net046 cn c VDD VSS net33 / TSINV pl=60n pw=340n nl=60n nw=240n
XI4 SI SE sen VDD VSS net046 / TSINV pl=60n pw=280n nl=60n nw=200n
XI3 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XI12 CK VDD VSS cn / INV pl=60n pw=340n nl=60n nw=240n
XI11 net25 VDD VSS net9 / INV pl=60n pw=340n nl=60n nw=240n
XI10 net25 VDD VSS Q / INV pl=60n pw=400n nl=60n nw=280n
XI9 cn VDD VSS c / INV pl=60n pw=340n nl=60n nw=240n
XI8 net33 VDD VSS net46 / INV pl=60n pw=340n nl=60n nw=240n
XI7 SE VDD VSS sen / INV pl=60n pw=340n nl=60n nw=240n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN0 Y B net15 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN2 net15 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP2 Y A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y B VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFTRQX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFTRQX3H7L CK D Q RN SE SI VDD VSS
*.PININFO CK:I D:I RN:I SE:I SI:I Q:O VDD:B VSS:B
XI3 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XI4 SI SE sen VDD VSS net046 / TSINV pl=60n pw=250n nl=60n nw=200n
XI5 net046 cn c VDD VSS net33 / TSINV pl=60n pw=360n nl=60n nw=260n
XI6 net9 cn c VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XI7 SE VDD VSS sen / INV pl=60n pw=340n nl=60n nw=240n
XI8 net33 VDD VSS net46 / INV pl=60n pw=360n nl=60n nw=260n
XI9 cn VDD VSS c / INV pl=60n pw=340n nl=60n nw=240n
XI10 net25 VDD VSS Q / INV pl=60n pw=600n nl=60n nw=420n
XI11 net25 VDD VSS net9 / INV pl=60n pw=360n nl=60n nw=260n
XI12 CK VDD VSS cn / INV pl=60n pw=340n nl=60n nw=240n
XI2 D RN VDD VSS net034 / NAND2 pl=60n pw=340n nl=60n nw=270n
XI0 c cn net46 net25 VDD VSS / TG pl=60n pw=360n nl=60n nw=260n
XI1 sen SE net034 net046 VDD VSS / TG pl=60n pw=360n nl=60n nw=260n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFX0P5H7L CK D Q QN SE SI VDD VSS
*.PININFO CK:I D:I SE:I SI:I Q:O QN:O VDD:B VSS:B
XXI14 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI18 SI SE sen VDD VSS net050 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI16 D sen SE VDD VSS net050 / TSINV pl=60n pw=300n nl=60n nw=220n
XXI9 net46 c cn VDD VSS net25 / TSINV pl=60n pw=280n nl=60n nw=200n
XXI15 net9 cn c VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI19 SE VDD VSS sen / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=280n nl=60n nw=200n
XXI13 cn VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net25 VDD VSS Q / INV pl=60n pw=280n nl=60n nw=200n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=280n nl=60n nw=200n
XXI5 net9 VDD VSS QN / INV pl=60n pw=280n nl=60n nw=200n
XXI4 CK VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
XXI17 cn c net050 net33 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFX1H7L CK D Q QN SE SI VDD VSS
*.PININFO CK:I D:I SE:I SI:I Q:O QN:O VDD:B VSS:B
XXI14 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI18 SI SE sen VDD VSS net050 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI16 D sen SE VDD VSS net050 / TSINV pl=60n pw=300n nl=60n nw=220n
XXI9 net46 c cn VDD VSS net25 / TSINV pl=60n pw=300n nl=60n nw=220n
XXI15 net9 cn c VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI19 SE VDD VSS sen / INV pl=60n pw=280n nl=60n nw=200n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=300n nl=60n nw=220n
XXI13 cn VDD VSS c / INV pl=60n pw=280n nl=60n nw=200n
XXI12 net25 VDD VSS Q / INV pl=60n pw=340n nl=60n nw=240n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=300n nl=60n nw=220n
XXI5 net9 VDD VSS QN / INV pl=60n pw=340n nl=60n nw=240n
XXI4 CK VDD VSS cn / INV pl=60n pw=280n nl=60n nw=200n
XXI17 cn c net050 net33 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFX2H7L CK D Q QN SE SI VDD VSS
*.PININFO CK:I D:I SE:I SI:I Q:O QN:O VDD:B VSS:B
XXI14 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI18 SI SE sen VDD VSS net050 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI16 D sen SE VDD VSS net050 / TSINV pl=60n pw=300n nl=60n nw=220n
XXI9 net46 c cn VDD VSS net25 / TSINV pl=60n pw=340n nl=60n nw=240n
XXI15 net9 cn c VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI19 SE VDD VSS sen / INV pl=60n pw=340n nl=60n nw=240n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=340n nl=60n nw=240n
XXI13 cn VDD VSS c / INV pl=60n pw=340n nl=60n nw=240n
XXI12 net25 VDD VSS Q / INV pl=60n pw=400n nl=60n nw=280n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=340n nl=60n nw=240n
XXI5 net9 VDD VSS QN / INV pl=60n pw=400n nl=60n nw=280n
XXI4 CK VDD VSS cn / INV pl=60n pw=340n nl=60n nw=240n
XXI17 cn c net050 net33 VDD VSS / TG pl=60n pw=300n nl=60n nw=220n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    SDFFX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT SDFFX3H7L CK D Q QN SE SI VDD VSS
*.PININFO CK:I D:I SE:I SI:I Q:O QN:O VDD:B VSS:B
XXI13 cn VDD VSS c / INV pl=60n pw=340n nl=60n nw=240n
XXI7 net33 VDD VSS net46 / INV pl=60n pw=360n nl=60n nw=260n
XXI12 net25 VDD VSS Q / INV pl=60n pw=600n nl=60n nw=420n
XXI19 SE VDD VSS sen / INV pl=60n pw=340n nl=60n nw=240n
XXI4 CK VDD VSS cn / INV pl=60n pw=340n nl=60n nw=240n
XXI5 net9 VDD VSS QN / INV pl=60n pw=600n nl=60n nw=420n
XXI10 net25 VDD VSS net9 / INV pl=60n pw=340n nl=60n nw=240n
XXI14 net46 c cn VDD VSS net33 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI18 SI SE sen VDD VSS net050 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI16 D sen SE VDD VSS net050 / TSINV pl=60n pw=340n nl=60n nw=240n
XXI9 net46 c cn VDD VSS net25 / TSINV pl=60n pw=360n nl=60n nw=260n
XXI15 net9 cn c VDD VSS net25 / TSINV pl=60n pw=150n nl=60n nw=150n
XXI17 cn c net050 net33 VDD VSS / TG pl=60n pw=340n nl=60n nw=240n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TBUFX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT TBUFX0P5H7L A OE VDD VSS Y
*.PININFO A:I OE:I Y:O VDD:B VSS:B
MNM0 net18 net39 VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MNM1 Y OE net18 VSS nm1p2_lvt_lp W=150n L=60n m=1
MPM0 Y OEN net17 VDD pm1p2_lvt_lp W=190n L=60n m=1
MPM1 net17 net39 VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XI2 OE VDD VSS OEN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XI1 A VDD VSS net39 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TBUFX0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT TBUFX0P7H7L A OE VDD VSS Y
*.PININFO A:I OE:I Y:O VDD:B VSS:B
MMNM0 net34 net39 VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN0 Y OE net34 VSS nm1p2_lvt_lp W=175n L=60n m=1
MMPM1 Y OEN net29 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM0 net29 net39 VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
XI1 OE VDD VSS OEN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI0 A VDD VSS net39 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TBUFX12H7L
* View Name:    schematic
************************************************************************

.SUBCKT TBUFX12H7L A OE VDD VSS Y
*.PININFO A:I OE:I Y:O VDD:B VSS:B
MNM0 net45 OEN VSS VSS nm1p2_lvt_lp W=1.74u L=60n m=1
MNM2 net45 A VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MNM1 Y net45 VSS VSS nm1p2_lvt_lp W=1.8u L=60n m=1
MPM0 Y net29 VDD VDD pm1p2_lvt_lp W=2.28u L=60n m=1
MPM1 net29 OE VDD VDD pm1p2_lvt_lp W=2.22u L=60n m=1
MPM2 net29 A VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
XI1 OE VDD VSS OEN / INV pl=6e-08 pw=7.6e-07 nl=6e-08 nw=6e-07
XI0 OE OEN net45 net29 VDD VSS / TG pl=6e-08 pw=7.6e-07 nl=6e-08 nw=6e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TBUFX16H7L
* View Name:    schematic
************************************************************************

.SUBCKT TBUFX16H7L A OE VDD VSS Y
*.PININFO A:I OE:I Y:O VDD:B VSS:B
MNM0 net45 OEN VSS VSS nm1p2_lvt_lp W=2.32u L=60n m=1
MNM2 net45 A VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MNM1 Y net45 VSS VSS nm1p2_lvt_lp W=2.4u L=60n m=1
MPM0 Y net29 VDD VDD pm1p2_lvt_lp W=3.04u L=60n m=1
MPM1 net29 OE VDD VDD pm1p2_lvt_lp W=2.96u L=60n m=1
MPM2 net29 A VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
XI1 OE VDD VSS OEN / INV pl=6e-08 pw=1.14e-06 nl=6e-08 nw=9e-07
XI0 OE OEN net45 net29 VDD VSS / TG pl=6e-08 pw=1.14e-06 nl=6e-08 nw=9e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TBUFX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT TBUFX1H7L A OE VDD VSS Y
*.PININFO A:I OE:I Y:O VDD:B VSS:B
MMNM0 net34 net39 VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN0 Y OE net34 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMPM1 Y OEN net29 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM0 net29 net39 VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
XI1 OE VDD VSS OEN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI0 A VDD VSS net39 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TBUFX1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT TBUFX1P4H7L A OE VDD VSS Y
*.PININFO A:I OE:I Y:O VDD:B VSS:B
MMNM0 net34 net39 VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN0 Y OE net34 VSS nm1p2_lvt_lp W=245n L=60n m=1
MMPM1 Y OEN net29 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM0 net29 net39 VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
XI1 OE VDD VSS OEN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI0 A VDD VSS net39 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TBUFX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT TBUFX2H7L A OE VDD VSS Y
*.PININFO A:I OE:I Y:O VDD:B VSS:B
MMNM0 net34 net39 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN0 Y OE net34 VSS nm1p2_lvt_lp W=300n L=60n m=1
MMPM1 Y OEN net29 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM0 net29 net39 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
XXI3 OE VDD VSS OEN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI0 A VDD VSS net39 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TBUFX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT TBUFX3H7L A OE VDD VSS Y
*.PININFO A:I OE:I Y:O VDD:B VSS:B
MNM2 net45 A VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MNM1 Y net45 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MNM0 net45 OEN VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MPM2 net29 A VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
MPM1 net29 OE VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MPM0 Y net29 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
XI1 OE VDD VSS OEN / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
XI0 OE OEN net45 net29 VDD VSS / TG pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TBUFX4H7L
* View Name:    schematic
************************************************************************

.SUBCKT TBUFX4H7L A OE VDD VSS Y
*.PININFO A:I OE:I Y:O VDD:B VSS:B
MNM2 net45 A VSS VSS nm1p2_lvt_lp W=250n L=60n m=1
MNM1 Y net45 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MNM0 net45 OEN VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MPM2 net29 A VDD VDD pm1p2_lvt_lp W=310n L=60n m=1
MPM1 net29 OE VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MPM0 Y net29 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
XI1 OE VDD VSS OEN / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
XI0 OE OEN net45 net29 VDD VSS / TG pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TBUFX6H7L
* View Name:    schematic
************************************************************************

.SUBCKT TBUFX6H7L A OE VDD VSS Y
*.PININFO A:I OE:I Y:O VDD:B VSS:B
MNM2 net45 A VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MNM1 Y net45 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MNM0 net45 OEN VSS VSS nm1p2_lvt_lp W=870n L=60n m=1
MPM2 net29 A VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MPM1 net29 OE VDD VDD pm1p2_lvt_lp W=1.11u L=60n m=1
MPM0 Y net29 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
XI0 OE OEN net45 net29 VDD VSS / TG pl=6e-08 pw=3.4e-07 nl=6e-08 nw=2.4e-07
XI1 OE VDD VSS OEN / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TBUFX8H7L
* View Name:    schematic
************************************************************************

.SUBCKT TBUFX8H7L A OE VDD VSS Y
*.PININFO A:I OE:I Y:O VDD:B VSS:B
XI1 OE VDD VSS OEN / INV pl=6e-08 pw=6.2e-07 nl=6e-08 nw=5e-07
XI0 OE OEN net45 net29 VDD VSS / TG pl=6e-08 pw=6.2e-07 nl=6e-08 nw=5e-07
MPM0 Y net29 VDD VDD pm1p2_lvt_lp W=1.52u L=60n m=1
MPM2 net29 A VDD VDD pm1p2_lvt_lp W=620n L=60n m=1
MPM1 net29 OE VDD VDD pm1p2_lvt_lp W=1.48u L=60n m=1
MNM2 net45 A VSS VSS nm1p2_lvt_lp W=500n L=60n m=1
MNM1 Y net45 VSS VSS nm1p2_lvt_lp W=1.2u L=60n m=1
MNM0 net45 OEN VSS VSS nm1p2_lvt_lp W=1.16u L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TIEHIH7L
* View Name:    schematic
************************************************************************

.SUBCKT TIELOH7L VDD VSS Z
*.PININFO Z:O VDD:B VSS:B
MMM1 Z net4 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMM0 net4 net4 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TIELOH7L
* View Name:    schematic
************************************************************************

.SUBCKT TIEHIH7L VDD VSS Z
*.PININFO Z:O VDD:B VSS:B
MMM0 Z net4 VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
MMM1 net4 net4 VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TINVX0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT TINVX0P5H7L A OE VDD VSS Y
*.PININFO A:I OE:I Y:O VDD:B VSS:B
MMNM0 net15 A VSS VSS nm1p2_lvt_lp W=150n L=60n m=1
MMN0 Y OE net15 VSS nm1p2_lvt_lp W=150n L=60n m=1
MMPM1 Y OEN net024 VDD pm1p2_lvt_lp W=190n L=60n m=1
MMPM0 net024 A VDD VDD pm1p2_lvt_lp W=190n L=60n m=1
XXI3 OE VDD VSS OEN / INV pl=6E-08 pw=1.9e-07 nl=6E-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TINVX0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT TINVX0P7H7L A OE VDD VSS Y
*.PININFO A:I OE:I Y:O VDD:B VSS:B
MNM0 net15 A VSS VSS nm1p2_lvt_lp W=175n L=60n m=1
MMN0 Y OE net15 VSS nm1p2_lvt_lp W=175n L=60n m=1
MPM0 Y OEN net024 VDD pm1p2_lvt_lp W=222n L=60n m=1
MMPM0 net024 A VDD VDD pm1p2_lvt_lp W=222n L=60n m=1
XXI3 OE VDD VSS OEN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TINVX12H7L
* View Name:    schematic
************************************************************************

.SUBCKT TINVX12H7L A OE VDD VSS Y
*.PININFO A:I OE:I Y:O VDD:B VSS:B
MNM0 net9 net27 VSS VSS nm1p2_lvt_lp W=1.8u L=60n m=1
MNM1 Y net9 VSS VSS nm1p2_lvt_lp W=1.8u L=60n m=1
MNM2 net9 OEN VSS VSS nm1p2_lvt_lp W=1.8u L=60n m=1
MPM2 Y net031 VDD VDD pm1p2_lvt_lp W=2.28u L=60n m=1
MPM1 net031 net27 VDD VDD pm1p2_lvt_lp W=2.28u L=60n m=1
MPM0 net031 OE VDD VDD pm1p2_lvt_lp W=2.28u L=60n m=1
XI2 OE VDD VSS OEN / INV pl=6E-08 pw=7.6e-07 nl=6E-08 nw=6e-07
XI1 A VDD VSS net27 / INV pl=6E-08 pw=2.28e-06 nl=6E-08 nw=1.8e-06
XI0 OE OEN net9 net031 VDD VSS / TG pl=6E-08 pw=2.22e-06 nl=6E-08 nw=1.74e-06
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TINVX16H7L
* View Name:    schematic
************************************************************************

.SUBCKT TINVX16H7L A OE VDD VSS Y
*.PININFO A:I OE:I Y:O VDD:B VSS:B
MNM0 net9 net27 VSS VSS nm1p2_lvt_lp W=2.4u L=60n m=1
MNM1 Y net9 VSS VSS nm1p2_lvt_lp W=2.4u L=60n m=1
MNM2 net9 OEN VSS VSS nm1p2_lvt_lp W=2.4u L=60n m=1
XI2 OE VDD VSS OEN / INV pl=6E-08 pw=1.14e-06 nl=6E-08 nw=9e-07
XI1 A VDD VSS net27 / INV pl=6E-08 pw=3.04e-06 nl=6E-08 nw=2.4e-06
MPM2 Y net031 VDD VDD pm1p2_lvt_lp W=3.04u L=60n m=1
MPM0 net031 OE VDD VDD pm1p2_lvt_lp W=3.04u L=60n m=1
MPM1 net031 net27 VDD VDD pm1p2_lvt_lp W=3.04u L=60n m=1
XI0 OE OEN net9 net031 VDD VSS / TG pl=6E-08 pw=2.96e-06 nl=6E-08 nw=2.32e-06
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TINVX1H7L
* View Name:    schematic
************************************************************************

.SUBCKT TINVX1H7L A OE VDD VSS Y
*.PININFO A:I OE:I Y:O VDD:B VSS:B
MMNM0 net15 A VSS VSS nm1p2_lvt_lp W=210n L=60n m=1
MMN0 Y OE net15 VSS nm1p2_lvt_lp W=210n L=60n m=1
MMPM1 Y OEN net024 VDD pm1p2_lvt_lp W=270n L=60n m=1
MMPM0 net024 A VDD VDD pm1p2_lvt_lp W=270n L=60n m=1
XXI3 OE VDD VSS OEN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TINVX1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT TINVX1P4H7L A OE VDD VSS Y
*.PININFO A:I OE:I Y:O VDD:B VSS:B
MNM0 net15 A VSS VSS nm1p2_lvt_lp W=245n L=60n m=1
MMN0 Y OE net15 VSS nm1p2_lvt_lp W=245n L=60n m=1
MPM0 Y OEN net024 VDD pm1p2_lvt_lp W=314n L=60n m=1
MMPM0 net024 A VDD VDD pm1p2_lvt_lp W=314n L=60n m=1
XXI3 OE VDD VSS OEN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TINVX2H7L
* View Name:    schematic
************************************************************************

.SUBCKT TINVX2H7L A OE VDD VSS Y
*.PININFO A:I OE:I Y:O VDD:B VSS:B
MNM0 net15 A VSS VSS nm1p2_lvt_lp W=300n L=60n m=1
MMN0 Y OE net15 VSS nm1p2_lvt_lp W=300n L=60n m=1
MPM0 Y OEN net024 VDD pm1p2_lvt_lp W=380n L=60n m=1
MMPM0 net024 A VDD VDD pm1p2_lvt_lp W=380n L=60n m=1
XXI3 OE VDD VSS OEN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TINVX3H7L
* View Name:    schematic
************************************************************************

.SUBCKT TINVX3H7L A OE VDD VSS Y
*.PININFO A:I OE:I Y:O VDD:B VSS:B
XI3 OE OEN net9 net031 VDD VSS / TG pl=6E-08 pw=5.7e-07 nl=6E-08 nw=4.5e-07
MNM7 net9 net27 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MNM9 Y net9 VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MNM8 net9 OEN VSS VSS nm1p2_lvt_lp W=450n L=60n m=1
MPM8 net031 OE VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MPM9 Y net031 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
MPM5 net031 net27 VDD VDD pm1p2_lvt_lp W=570n L=60n m=1
XI5 OE VDD VSS OEN / INV pl=6E-08 pw=3.1e-07 nl=6E-08 nw=2.5e-07
XI4 A VDD VSS net27 / INV pl=6E-08 pw=5.7e-07 nl=6E-08 nw=4.5e-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TINVX4H7L
* View Name:    schematic
************************************************************************

.SUBCKT TINVX4H7L A OE VDD VSS Y
*.PININFO A:I OE:I Y:O VDD:B VSS:B
XI3 OE OEN net9 net031 VDD VSS / TG pl=6E-08 pw=7.6e-07 nl=6E-08 nw=6e-07
MNM7 net9 net27 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MNM6 net9 OEN VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MNM5 Y net9 VSS VSS nm1p2_lvt_lp W=600n L=60n m=1
MPM7 Y net031 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MPM6 net031 OE VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
MPM5 net031 net27 VDD VDD pm1p2_lvt_lp W=760n L=60n m=1
XI5 OE VDD VSS OEN / INV pl=6E-08 pw=3.1e-07 nl=6E-08 nw=2.5e-07
XI4 A VDD VSS net27 / INV pl=6E-08 pw=7.6e-07 nl=6E-08 nw=6e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TINVX6H7L
* View Name:    schematic
************************************************************************

.SUBCKT TINVX6H7L A OE VDD VSS Y
*.PININFO A:I OE:I Y:O VDD:B VSS:B
MNM7 Y net9 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MNM6 net9 OEN VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MNM5 net9 net27 VSS VSS nm1p2_lvt_lp W=900n L=60n m=1
MPM7 Y net031 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MPM6 net031 OE VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
MPM5 net031 net27 VDD VDD pm1p2_lvt_lp W=1.14u L=60n m=1
XI5 A VDD VSS net27 / INV pl=6E-08 pw=1.14e-06 nl=6E-08 nw=9e-07
XI3 OE VDD VSS OEN / INV pl=6E-08 pw=3.8e-07 nl=6E-08 nw=3e-07
XI4 OE OEN net9 net031 VDD VSS / TG pl=6E-08 pw=1.14e-06 nl=6E-08 nw=9e-07
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    TINVX8H7L
* View Name:    schematic
************************************************************************

.SUBCKT TINVX8H7L A OE VDD VSS Y
*.PININFO A:I OE:I Y:O VDD:B VSS:B
MPM0 net031 OE VDD VDD pm1p2_lvt_lp W=1.52u L=60n m=1
MMPM0 Y net031 VDD VDD pm1p2_lvt_lp W=1.52u L=60n m=1
MPM1 net031 net27 VDD VDD pm1p2_lvt_lp W=1.52u L=60n m=1
MNM2 net9 OEN VSS VSS nm1p2_lvt_lp W=1.2u L=60n m=1
MNM0 net9 net27 VSS VSS nm1p2_lvt_lp W=1.2u L=60n m=1
MNM1 Y net9 VSS VSS nm1p2_lvt_lp W=1.2u L=60n m=1
XXI3 OE VDD VSS OEN / INV pl=6E-08 pw=6.2e-07 nl=6E-08 nw=5e-07
XXI7 A VDD VSS net27 / INV pl=6E-08 pw=1.52e-06 nl=6E-08 nw=1.2e-06
XXI6 OE OEN net9 net031 VDD VSS / TG pl=6E-08 pw=1.48e-06 nl=6E-08 nw=1.16e-06
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XNOR2X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT XNOR2X0P5H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
XXI4 A AN BN net19 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI9 net19 VDD VSS Y / INV pl=60n pw=190n nl=60n nw=150n
XXI7 B VDD VSS BN / INV pl=60n pw=190n nl=60n nw=150n
XXI0 A VDD VSS AN / INV pl=60n pw=190n nl=60n nw=150n
XXI10 BN AN A VDD VSS net19 / TSINV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XNOR2X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT XNOR2X0P7H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
XXI4 A AN BN net19 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI0 A VDD VSS AN / INV pl=60n pw=190n nl=60n nw=150n
XXI7 B VDD VSS BN / INV pl=60n pw=190n nl=60n nw=150n
XXI9 net19 VDD VSS Y / INV pl=60n pw=222n nl=60n nw=174n
XXI10 BN AN A VDD VSS net19 / TSINV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XNOR2X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT XNOR2X1H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
XXI4 A AN BN net19 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI9 net19 VDD VSS Y / INV pl=60n pw=270n nl=60n nw=210n
XXI7 B VDD VSS BN / INV pl=60n pw=190n nl=60n nw=150n
XXI0 A VDD VSS AN / INV pl=60n pw=190n nl=60n nw=150n
XXI10 BN AN A VDD VSS net19 / TSINV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XNOR2X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT XNOR2X1P4H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
XXI4 A AN BN net19 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI0 A VDD VSS AN / INV pl=60n pw=190n nl=60n nw=150n
XXI7 B VDD VSS BN / INV pl=60n pw=190n nl=60n nw=150n
XXI9 net19 VDD VSS Y / INV pl=60n pw=314n nl=60n nw=246n
XXI10 BN AN A VDD VSS net19 / TSINV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XNOR2X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT XNOR2X2H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
XXI4 A AN BN net19 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI0 A VDD VSS AN / INV pl=60n pw=190n nl=60n nw=150n
XXI7 B VDD VSS BN / INV pl=60n pw=190n nl=60n nw=150n
XXI9 net19 VDD VSS Y / INV pl=60n pw=380n nl=60n nw=300n
XXI10 BN AN A VDD VSS net19 / TSINV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XNOR2X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT XNOR2X3H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
XXI4 A AN BN net19 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI0 A VDD VSS AN / INV pl=60n pw=200n nl=60n nw=160n
XXI7 B VDD VSS BN / INV pl=60n pw=250n nl=60n nw=200n
XXI9 net19 VDD VSS Y / INV pl=60n pw=570n nl=60n nw=450n
XXI10 BN AN A VDD VSS net19 / TSINV pl=60n pw=250n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XNOR2X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT XNOR2X4H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
XXI10 BN AN A VDD VSS net19 / TSINV pl=60n pw=310n nl=60n nw=250n
XXI9 net19 VDD VSS Y / INV pl=60n pw=760n nl=60n nw=600n
XXI7 B VDD VSS BN / INV pl=60n pw=310n nl=60n nw=250n
XXI0 A VDD VSS AN / INV pl=60n pw=210n nl=60n nw=170n
XXI4 A AN BN net19 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XNOR2X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT XNOR2X6H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
XXI4 A AN BN net19 VDD VSS / TG pl=60n pw=210n nl=60n nw=170n
XXI0 A VDD VSS AN / INV pl=60n pw=250n nl=60n nw=200n
XXI7 B VDD VSS BN / INV pl=60n pw=380n nl=60n nw=300n
XXI9 net19 VDD VSS Y / INV pl=60n pw=1140n nl=60n nw=900n
XXI10 BN AN A VDD VSS net19 / TSINV pl=60n pw=310n nl=60n nw=250n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XNOR3X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT XNOR3X0P5H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
XXI16 AN A BN net45 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI14 net57 net45 CN net49 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI18 BN A AN VDD VSS net45 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI13 CN net45 net57 VDD VSS net49 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI15 net45 VDD VSS net57 / INV pl=60n pw=190n nl=60n nw=150n
XXI17 B VDD VSS BN / INV pl=60n pw=190n nl=60n nw=150n
XXI11 net49 VDD VSS Y / INV pl=60n pw=190n nl=60n nw=150n
XXI19 A VDD VSS AN / INV pl=60n pw=190n nl=60n nw=150n
XXI12 C VDD VSS CN / INV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XNOR3X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT XNOR3X0P7H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
XXI16 AN A BN net45 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI14 net57 net45 CN net49 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI18 BN A AN VDD VSS net45 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI13 CN net45 net57 VDD VSS net49 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI15 net45 VDD VSS net57 / INV pl=60n pw=190n nl=60n nw=150n
XXI17 B VDD VSS BN / INV pl=60n pw=190n nl=60n nw=150n
XXI11 net49 VDD VSS Y / INV pl=60n pw=222n nl=60n nw=174n
XXI19 A VDD VSS AN / INV pl=60n pw=190n nl=60n nw=150n
XXI12 C VDD VSS CN / INV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XNOR3X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT XNOR3X1H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
XXI16 AN A BN net45 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI14 net57 net45 CN net49 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI18 BN A AN VDD VSS net45 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI13 CN net45 net57 VDD VSS net49 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI15 net45 VDD VSS net57 / INV pl=60n pw=190n nl=60n nw=150n
XXI17 B VDD VSS BN / INV pl=60n pw=190n nl=60n nw=150n
XXI11 net49 VDD VSS Y / INV pl=60n pw=270n nl=60n nw=210n
XXI19 A VDD VSS AN / INV pl=60n pw=190n nl=60n nw=150n
XXI12 C VDD VSS CN / INV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XNOR3X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT XNOR3X1P4H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
XXI16 AN A BN net45 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI14 net57 net45 CN net49 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI18 BN A AN VDD VSS net45 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI13 CN net45 net57 VDD VSS net49 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI15 net45 VDD VSS net57 / INV pl=60n pw=190n nl=60n nw=150n
XXI17 B VDD VSS BN / INV pl=60n pw=220n nl=60n nw=175n
XXI11 net49 VDD VSS Y / INV pl=60n pw=325n nl=60n nw=255n
XXI19 A VDD VSS AN / INV pl=60n pw=190n nl=60n nw=150n
XXI12 C VDD VSS CN / INV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XNOR3X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT XNOR3X2H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
XXI16 AN A BN net45 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI14 net57 net45 CN net49 VDD VSS / TG pl=60n pw=190n nl=60n nw=150n
XXI18 BN A AN VDD VSS net45 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI13 CN net45 net57 VDD VSS net49 / TSINV pl=60n pw=190n nl=60n nw=150n
XXI15 net45 VDD VSS net57 / INV pl=60n pw=190n nl=60n nw=150n
XXI17 B VDD VSS BN / INV pl=60n pw=250n nl=60n nw=200n
XXI11 net49 VDD VSS Y / INV pl=60n pw=380n nl=60n nw=300n
XXI19 A VDD VSS AN / INV pl=60n pw=190n nl=60n nw=150n
XXI12 C VDD VSS CN / INV pl=60n pw=190n nl=60n nw=150n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XNOR3X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT XNOR3X3H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
XXI16 AN A BN net45 VDD VSS / TG pl=60n pw=220n nl=60n nw=175n
XXI14 net57 net45 CN net49 VDD VSS / TG pl=60n pw=220n nl=60n nw=175n
XXI18 BN A AN VDD VSS net45 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI13 CN net45 net57 VDD VSS net49 / TSINV pl=60n pw=250n nl=60n nw=200n
XXI15 net45 VDD VSS net57 / INV pl=60n pw=250n nl=60n nw=200n
XXI17 B VDD VSS BN / INV pl=60n pw=280n nl=60n nw=225n
XXI11 net49 VDD VSS Y / INV pl=60n pw=570n nl=60n nw=450n
XXI19 A VDD VSS AN / INV pl=60n pw=250n nl=60n nw=200n
XXI12 C VDD VSS CN / INV pl=60n pw=250n nl=60n nw=200n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XNOR3X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT XNOR3X4H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
XXI15 net45 VDD VSS net57 / INV pl=60n pw=310n nl=60n nw=250n
XXI17 B VDD VSS BN / INV pl=60n pw=310n nl=60n nw=250n
XXI12 C VDD VSS CN / INV pl=60n pw=310n nl=60n nw=250n
XXI19 A VDD VSS AN / INV pl=60n pw=310n nl=60n nw=250n
XXI11 net49 VDD VSS Y / INV pl=60n pw=760n nl=60n nw=600n
XXI13 CN net45 net57 VDD VSS net49 / TSINV pl=60n pw=310n nl=60n nw=250n
XXI18 BN A AN VDD VSS net45 / TSINV pl=60n pw=310n nl=60n nw=250n
XXI14 net57 net45 CN net49 VDD VSS / TG pl=60n pw=250n nl=60n nw=200n
XXI16 AN A BN net45 VDD VSS / TG pl=60n pw=250n nl=60n nw=200n
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XNOR3X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT XNOR3X6H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
XXI11 net49 VDD VSS Y / INV pl=60n pw=1140n nl=60n nw=900n
XXI19 A VDD VSS AN / INV pl=60n pw=310n nl=60n nw=250n
XXI12 C VDD VSS CN / INV pl=60n pw=310n nl=60n nw=250n
XXI17 B VDD VSS BN / INV pl=60n pw=310n nl=60n nw=250n
XXI15 net45 VDD VSS net57 / INV pl=60n pw=310n nl=60n nw=250n
XXI18 BN A AN VDD VSS net45 / TSINV pl=60n pw=310n nl=60n nw=250n
XXI13 CN net45 net57 VDD VSS net49 / TSINV pl=60n pw=310n nl=60n nw=250n
XXI16 AN A BN net45 VDD VSS / TG pl=60n pw=250n nl=60n nw=200n
XXI14 net57 net45 CN net49 VDD VSS / TG pl=60n pw=250n nl=60n nw=200n
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XOR2X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT XOR2X0P5H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
XI0 AN A BN net19 VDD VSS / TG pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XI6 net19 VDD VSS Y / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XI1 B VDD VSS BN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XI4 A VDD VSS AN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XI3 BN A AN VDD VSS net19 / TSINV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XOR2X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT XOR2X0P7H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
XI0 AN A BN net19 VDD VSS / TG pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XI6 net19 VDD VSS Y / INV pl=6e-08 pw=2.22e-07 nl=6e-08 nw=1.74e-07
XI1 B VDD VSS BN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XI4 A VDD VSS AN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XI3 BN A AN VDD VSS net19 / TSINV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XOR2X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT XOR2X1H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
XI0 AN A BN net19 VDD VSS / TG pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XI5 net19 VDD VSS Y / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
XI1 B VDD VSS BN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XI4 A VDD VSS AN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XI3 BN A AN VDD VSS net19 / TSINV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XOR2X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT XOR2X1P4H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
XI0 AN A BN net19 VDD VSS / TG pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XI5 net19 VDD VSS Y / INV pl=6e-08 pw=3.14e-07 nl=6e-08 nw=2.46e-07
XI1 B VDD VSS BN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XI4 A VDD VSS AN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XI3 BN A AN VDD VSS net19 / TSINV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XOR2X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT XOR2X2H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
XI0 AN A BN net19 VDD VSS / TG pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XI1 B VDD VSS BN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XI4 A VDD VSS AN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XI2 net19 VDD VSS Y / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
XI3 BN A AN VDD VSS net19 / TSINV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XOR2X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT XOR2X3H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
XI0 AN A BN net19 VDD VSS / TG pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XI1 B VDD VSS BN / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
XI4 A VDD VSS AN / INV pl=6e-08 pw=2.1e-07 nl=6e-08 nw=1.7e-07
XI2 net19 VDD VSS Y / INV pl=6e-08 pw=5.7e-07 nl=6e-08 nw=4.5e-07
XI3 BN A AN VDD VSS net19 / TSINV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XOR2X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT XOR2X4H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
XI0 AN A BN net19 VDD VSS / TG pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XI1 B VDD VSS BN / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
XI4 A VDD VSS AN / INV pl=6e-08 pw=2.1e-07 nl=6e-08 nw=1.7e-07
XI2 net19 VDD VSS Y / INV pl=6e-08 pw=7.6e-07 nl=6e-08 nw=6e-07
XI3 BN A AN VDD VSS net19 / TSINV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XOR2X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT XOR2X6H7L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
XI0 AN A BN net19 VDD VSS / TG pl=6e-08 pw=2.1e-07 nl=6e-08 nw=1.7e-07
XI2 net19 VDD VSS Y / INV pl=6e-08 pw=11.4e-07 nl=6e-08 nw=9e-07
XI1 B VDD VSS BN / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
XI4 A VDD VSS AN / INV pl=6e-08 pw=2.5e-07 nl=6e-08 nw=2e-07
XI3 BN A AN VDD VSS net19 / TSINV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XOR3X0P5H7L
* View Name:    schematic
************************************************************************

.SUBCKT XOR3X0P5H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
XXI16 A AN net55 net45 VDD VSS / TG pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI14 net57 net45 net59 net49 VDD VSS / TG pl=6e-08 pw=1.9e-07 nl=6e-08
+ nw=1.5e-07
XXI15 net45 VDD VSS net57 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI17 B VDD VSS net55 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XI0 net49 VDD VSS Y / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI19 A VDD VSS AN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI12 C VDD VSS net59 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI18 net55 AN A VDD VSS net45 / TSINV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI13 net59 net45 net57 VDD VSS net49 / TSINV pl=6e-08 pw=1.9e-07 nl=6e-08
+ nw=1.5e-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XOR3X0P7H7L
* View Name:    schematic
************************************************************************

.SUBCKT XOR3X0P7H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
XXI16 A AN net55 net45 VDD VSS / TG pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI14 net57 net45 net59 net49 VDD VSS / TG pl=6e-08 pw=1.9e-07 nl=6e-08
+ nw=1.5e-07
XXI15 net45 VDD VSS net57 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI17 B VDD VSS net55 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI11 net49 VDD VSS Y / INV pl=6e-08 pw=2.22e-07 nl=6e-08 nw=1.74e-07
XXI19 A VDD VSS AN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI12 C VDD VSS net59 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI18 net55 AN A VDD VSS net45 / TSINV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI13 net59 net45 net57 VDD VSS net49 / TSINV pl=6e-08 pw=1.9e-07 nl=6e-08
+ nw=1.5e-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XOR3X1H7L
* View Name:    schematic
************************************************************************

.SUBCKT XOR3X1H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
XXI16 A AN net55 net45 VDD VSS / TG pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI14 net57 net45 net59 net49 VDD VSS / TG pl=6e-08 pw=1.9e-07 nl=6e-08
+ nw=1.5e-07
XXI15 net45 VDD VSS net57 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI17 B VDD VSS net55 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI11 net49 VDD VSS Y / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
XXI19 A VDD VSS AN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI12 C VDD VSS net59 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI18 net55 AN A VDD VSS net45 / TSINV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI13 net59 net45 net57 VDD VSS net49 / TSINV pl=6e-08 pw=1.9e-07 nl=6e-08
+ nw=1.5e-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XOR3X1P4H7L
* View Name:    schematic
************************************************************************

.SUBCKT XOR3X1P4H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
XXI16 A AN net55 net45 VDD VSS / TG pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI14 net57 net45 net59 net49 VDD VSS / TG pl=6e-08 pw=1.9e-07 nl=6e-08
+ nw=1.5e-07
XXI15 net45 VDD VSS net57 / INV pl=6e-08 pw=2.1e-07 nl=6e-08 nw=1.7e-07
XXI17 B VDD VSS net55 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI11 net49 VDD VSS Y / INV pl=6e-08 pw=3.14e-07 nl=6e-08 nw=2.46e-07
XXI19 A VDD VSS AN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI12 C VDD VSS net59 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI18 net55 AN A VDD VSS net45 / TSINV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI13 net59 net45 net57 VDD VSS net49 / TSINV pl=6e-08 pw=1.9e-07 nl=6e-08
+ nw=1.5e-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XOR3X2H7L
* View Name:    schematic
************************************************************************

.SUBCKT XOR3X2H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
XXI16 A AN net55 net45 VDD VSS / TG pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI14 net57 net45 net59 net49 VDD VSS / TG pl=6e-08 pw=1.9e-07 nl=6e-08
+ nw=1.5e-07
XXI15 net45 VDD VSS net57 / INV pl=6e-08 pw=2.5e-07 nl=6e-08 nw=2e-07
XXI17 B VDD VSS net55 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI11 net49 VDD VSS Y / INV pl=6e-08 pw=3.8e-07 nl=6e-08 nw=3e-07
XXI19 A VDD VSS AN / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI12 C VDD VSS net59 / INV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI18 net55 AN A VDD VSS net45 / TSINV pl=6e-08 pw=1.9e-07 nl=6e-08 nw=1.5e-07
XXI13 net59 net45 net57 VDD VSS net49 / TSINV pl=6e-08 pw=1.9e-07 nl=6e-08
+ nw=1.5e-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XOR3X3H7L
* View Name:    schematic
************************************************************************

.SUBCKT XOR3X3H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
XXI16 A AN net55 net45 VDD VSS / TG pl=6e-08 pw=2.1e-07 nl=6e-08 nw=1.7e-07
XXI14 net57 net45 net59 net49 VDD VSS / TG pl=6e-08 pw=2.1e-07 nl=6e-08
+ nw=1.7e-07
XXI15 net45 VDD VSS net57 / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
XI0 B VDD VSS net55 / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
XXI11 net49 VDD VSS Y / INV pl=6e-08 pw=5.7e-07 nl=6e-08 nw=4.5e-07
XI1 A VDD VSS AN / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
XI2 C VDD VSS net59 / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
XXI18 net55 AN A VDD VSS net45 / TSINV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
XI3 net59 net45 net57 VDD VSS net49 / TSINV pl=6e-08 pw=2.7e-07 nl=6e-08
+ nw=2.1e-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XOR3X4H7L
* View Name:    schematic
************************************************************************

.SUBCKT XOR3X4H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
XXI16 A AN net55 net45 VDD VSS / TG pl=6e-08 pw=2.5e-07 nl=6e-08 nw=1.9e-07
XXI14 net57 net45 net59 net49 VDD VSS / TG pl=6e-08 pw=2.5e-07 nl=6e-08
+ nw=2e-07
XXI15 net45 VDD VSS net57 / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
XXI17 B VDD VSS net55 / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
XXI11 net49 VDD VSS Y / INV pl=6e-08 pw=7.6e-07 nl=6e-08 nw=6e-07
XXI19 A VDD VSS AN / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
XXI12 C VDD VSS net59 / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
XXI18 net55 AN A VDD VSS net45 / TSINV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
XXI13 net59 net45 net57 VDD VSS net49 / TSINV pl=6e-08 pw=3.1e-07 nl=6e-08
+ nw=2.5e-07
.ENDS

************************************************************************
* Library Name: ICSCORE
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG CK CKN D Q VDD VSS
*.PININFO CK:I CKN:I D:B Q:B VDD:B VSS:B
MMN0 D CK Q VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP0 D CKN Q VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************

************************************************************************



************************************************************************
* Library Name: ICSCORE
* Cell Name:    TSINV
* View Name:    schematic
************************************************************************

.SUBCKT TSINV A CK CKN VDD VSS Y
*.PININFO A:I CK:I CKN:I VDD:B VSS:B Y:B
MMN0 Y CK net18 VSS nm1p2_lvt_lp W=nw L=nl m=1
MMN1 net18 A VSS VSS nm1p2_lvt_lp W=nw L=nl m=1
MMP1 net024 A VDD VDD pm1p2_lvt_lp W=pw L=pl m=1
MMP0 Y CKN net024 VDD pm1p2_lvt_lp W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: ICSN55H7LVT
* Cell Name:    XOR3X6H7L
* View Name:    schematic
************************************************************************

.SUBCKT XOR3X6H7L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
XXI16 A AN net55 net45 VDD VSS / TG pl=6e-08 pw=2.5e-07 nl=6e-08 nw=1.9e-07
XXI14 net57 net45 net59 net49 VDD VSS / TG pl=6e-08 pw=2.5e-07 nl=6e-08
+ nw=2e-07
XXI15 net45 VDD VSS net57 / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
XXI17 B VDD VSS net55 / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
XXI11 net49 VDD VSS Y / INV pl=6e-08 pw=11.4e-07 nl=6e-08 nw=9e-07
XXI19 A VDD VSS AN / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
XXI12 C VDD VSS net59 / INV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
XXI18 net55 AN A VDD VSS net45 / TSINV pl=6e-08 pw=3.1e-07 nl=6e-08 nw=2.5e-07
XXI13 net59 net45 net57 VDD VSS net49 / TSINV pl=6e-08 pw=3.1e-07 nl=6e-08
+ nw=2.5e-07
.ENDS
.SUBCKT ANT2H7L VSS VDD A
** N=3 EP=3 IP=0 FDC=3
D0 VSS A dio_1p2_np_pw_lvt_lp AREA=8.7e-14 PJ=1.18e-06 m=1 l=3e-07 w=2.9e-07 $X=55 $Y=155 $D=163
D1 A VDD dio_1p2_pp_nw_lvt_lp AREA=1.1e-13 PJ=1.35e-06 m=1 l=4e-07 w=2.75e-07 $X=55 $Y=775 $D=164
.ENDS

.SUBCKT ANT4H7L VSS VDD A
** N=3 EP=3 IP=0 FDC=3
D0 VSS A dio_1p2_np_pw_lvt_lp AREA=2.07e-13 PJ=1.98e-06 m=1 l=6.9e-07 w=3e-07 $X=55 $Y=165 $D=163
D1 A VDD dio_1p2_pp_nw_lvt_lp AREA=2.622e-13 PJ=2.074e-06 m=1 l=6e-07 w=4.37e-07 $X=55 $Y=765 $D=164
.ENDS
