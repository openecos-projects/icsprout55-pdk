# Copyright 2025 ICsprout Integrated Circuit Co., Ltd.
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO ADDFX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFX1H7R 0 0 ;
  SIZE 4.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.8 1.48 ;
        RECT 4.215 1.19 4.355 1.48 ;
        RECT 3.71 1.19 3.8 1.48 ;
        RECT 1.825 1.085 1.915 1.48 ;
        RECT 0.07 0.855 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.8 0.08 ;
        RECT 4.24 -0.08 4.33 0.375 ;
        RECT 3.7 -0.08 3.79 0.36 ;
        RECT 1.81 -0.08 1.9 0.33 ;
        RECT 0.045 -0.08 0.185 0.32 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.555 0.545 0.78 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.425 0.175 0.65 ;
      LAYER MET2 ;
        RECT 0.05 0.23 0.15 0.76 ;
      LAYER VIA1 ;
        RECT 0.055 0.455 0.145 0.545 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.663 0.53 3.02 0.62 ;
        RECT 2.558 0.511 2.701 0.534 ;
        RECT 1.56 0.481 2.663 0.515 ;
        RECT 2.642 0.53 3.02 0.61 ;
        RECT 1.56 0.448 2.642 0.515 ;
        RECT 2.596 0.53 3.02 0.576 ;
        RECT 1.56 0.425 2.596 0.515 ;
        RECT 2.025 0.425 2.285 0.56 ;
      LAYER MET2 ;
        RECT 2.05 0.23 2.15 0.76 ;
      LAYER VIA1 ;
        RECT 2.055 0.455 2.145 0.545 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.975 0.225 4.145 0.375 ;
        RECT 3.975 0.225 4.065 0.92 ;
      LAYER MET2 ;
        RECT 4.05 0.18 4.15 0.56 ;
      LAYER VIA1 ;
        RECT 4.055 0.255 4.145 0.345 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.505 0.255 4.595 0.935 ;
        RECT 4.425 0.255 4.595 0.345 ;
      LAYER MET2 ;
        RECT 4.45 0.18 4.55 0.56 ;
      LAYER VIA1 ;
        RECT 4.455 0.255 4.545 0.345 ;
    END
  END S
  OBS
    LAYER MET1 ;
      RECT 3.795 1.01 4.415 1.1 ;
      RECT 4.325 0.585 4.415 1.1 ;
      RECT 3.795 0.54 3.885 1.1 ;
      RECT 2.49 0.82 2.63 0.91 ;
      RECT 2.49 0.82 2.632 0.909 ;
      RECT 2.49 0.82 2.67 0.889 ;
      RECT 3.16 0.35 3.25 0.87 ;
      RECT 2.592 0.801 3.25 0.87 ;
      RECT 2.632 0.78 3.25 0.87 ;
      RECT 2.63 0.781 3.25 0.87 ;
      RECT 3.16 0.54 3.885 0.63 ;
      RECT 2.739 0.35 3.25 0.44 ;
      RECT 2.718 0.301 2.739 0.43 ;
      RECT 2.672 0.268 2.718 0.396 ;
      RECT 2.634 0.331 2.777 0.354 ;
      RECT 2.49 0.245 2.672 0.335 ;
      RECT 2.005 1.14 3.61 1.23 ;
      RECT 2.005 0.905 2.095 1.23 ;
      RECT 0.635 1.035 1.735 1.125 ;
      RECT 1.645 0.905 1.735 1.125 ;
      RECT 0.635 0.395 0.725 1.125 ;
      RECT 1.645 0.905 2.095 0.995 ;
      RECT 0.505 0.895 0.725 0.985 ;
      RECT 0.635 0.395 1.32 0.485 ;
      RECT 1.18 0.36 1.32 0.485 ;
      RECT 0.62 0.336 0.635 0.465 ;
      RECT 0.576 0.392 0.686 0.435 ;
      RECT 0.576 0.367 0.681 0.435 ;
      RECT 0.53 0.19 0.62 0.39 ;
      RECT 3.43 0.17 3.52 0.36 ;
      RECT 2.815 0.17 3.52 0.26 ;
      RECT 2.8 0.96 3.52 1.05 ;
      RECT 3.43 0.85 3.52 1.05 ;
      RECT 1.62 0.65 2.379 0.74 ;
      RECT 1.595 0.65 2.381 0.728 ;
      RECT 1.595 0.65 2.419 0.719 ;
      RECT 0.845 0.625 1.633 0.715 ;
      RECT 2.381 0.61 2.525 0.7 ;
      RECT 2.341 0.631 2.525 0.7 ;
      RECT 2.379 0.611 2.381 0.739 ;
      RECT 0.845 0.637 1.658 0.715 ;
      RECT 0.845 0.575 0.935 0.715 ;
      RECT 0.755 0.17 0.9 0.305 ;
      RECT 0.755 0.17 1.57 0.26 ;
      RECT 0.885 0.855 1.555 0.945 ;
      RECT 1.465 0.805 1.555 0.945 ;
  END
END ADDFX1H7R

MACRO ADDFX1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFX1P4H7R 0 0 ;
  SIZE 4.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.8 1.48 ;
        RECT 4.215 1.19 4.355 1.48 ;
        RECT 3.71 1.19 3.8 1.48 ;
        RECT 1.82 1.085 1.91 1.48 ;
        RECT 0.07 0.855 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.8 0.08 ;
        RECT 4.24 -0.08 4.33 0.345 ;
        RECT 3.7 -0.08 3.79 0.33 ;
        RECT 1.805 -0.08 1.895 0.33 ;
        RECT 0.045 -0.08 0.185 0.32 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.555 0.545 0.78 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.425 0.175 0.65 ;
      LAYER MET2 ;
        RECT 0.05 0.23 0.15 0.76 ;
      LAYER VIA1 ;
        RECT 0.055 0.455 0.145 0.545 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.658 0.53 3.02 0.62 ;
        RECT 2.553 0.511 2.696 0.534 ;
        RECT 1.555 0.481 2.658 0.515 ;
        RECT 2.637 0.53 3.02 0.61 ;
        RECT 1.555 0.448 2.637 0.515 ;
        RECT 2.591 0.53 3.02 0.576 ;
        RECT 1.555 0.425 2.591 0.515 ;
        RECT 2.02 0.425 2.28 0.56 ;
      LAYER MET2 ;
        RECT 2.05 0.23 2.15 0.76 ;
      LAYER VIA1 ;
        RECT 2.055 0.455 2.145 0.545 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.05 0.225 4.145 0.375 ;
        RECT 3.975 0.285 4.065 0.92 ;
      LAYER MET2 ;
        RECT 4.05 0.18 4.15 0.56 ;
      LAYER VIA1 ;
        RECT 4.055 0.255 4.145 0.345 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.505 0.255 4.595 0.935 ;
        RECT 4.425 0.255 4.595 0.345 ;
      LAYER MET2 ;
        RECT 4.45 0.18 4.55 0.56 ;
      LAYER VIA1 ;
        RECT 4.455 0.255 4.545 0.345 ;
    END
  END S
  OBS
    LAYER MET1 ;
      RECT 3.795 1.01 4.415 1.1 ;
      RECT 4.325 0.585 4.415 1.1 ;
      RECT 3.795 0.54 3.885 1.1 ;
      RECT 2.485 0.82 2.625 0.91 ;
      RECT 2.485 0.82 2.627 0.909 ;
      RECT 2.485 0.82 2.665 0.889 ;
      RECT 3.16 0.35 3.25 0.87 ;
      RECT 2.587 0.801 3.25 0.87 ;
      RECT 2.627 0.78 3.25 0.87 ;
      RECT 2.625 0.781 3.25 0.87 ;
      RECT 3.16 0.54 3.885 0.63 ;
      RECT 2.734 0.35 3.25 0.44 ;
      RECT 2.713 0.301 2.734 0.43 ;
      RECT 2.667 0.268 2.713 0.396 ;
      RECT 2.629 0.331 2.772 0.354 ;
      RECT 2.485 0.245 2.667 0.335 ;
      RECT 2 1.14 3.61 1.23 ;
      RECT 2 0.905 2.09 1.23 ;
      RECT 0.635 1.035 1.73 1.125 ;
      RECT 1.64 0.905 1.73 1.125 ;
      RECT 0.635 0.395 0.725 1.125 ;
      RECT 1.64 0.905 2.09 0.995 ;
      RECT 0.505 0.895 0.725 0.985 ;
      RECT 0.635 0.395 1.315 0.485 ;
      RECT 1.175 0.36 1.315 0.485 ;
      RECT 0.62 0.336 0.635 0.465 ;
      RECT 0.576 0.392 0.686 0.435 ;
      RECT 0.576 0.367 0.681 0.435 ;
      RECT 0.53 0.19 0.62 0.39 ;
      RECT 3.43 0.17 3.52 0.33 ;
      RECT 2.815 0.17 3.52 0.26 ;
      RECT 2.8 0.96 3.52 1.05 ;
      RECT 3.43 0.85 3.52 1.05 ;
      RECT 1.618 0.65 2.374 0.74 ;
      RECT 1.593 0.65 2.376 0.728 ;
      RECT 1.593 0.65 2.414 0.719 ;
      RECT 0.84 0.625 1.631 0.715 ;
      RECT 2.376 0.61 2.52 0.7 ;
      RECT 2.336 0.631 2.52 0.7 ;
      RECT 2.374 0.611 2.376 0.739 ;
      RECT 0.84 0.637 1.656 0.715 ;
      RECT 0.84 0.575 0.93 0.715 ;
      RECT 0.755 0.17 0.9 0.305 ;
      RECT 0.755 0.17 1.565 0.26 ;
      RECT 0.88 0.855 1.55 0.945 ;
      RECT 1.46 0.805 1.55 0.945 ;
  END
END ADDFX1P4H7R

MACRO ADDFX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFX2H7R 0 0 ;
  SIZE 5 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5 1.48 ;
        RECT 4.755 0.835 4.845 1.48 ;
        RECT 4.215 1.19 4.355 1.48 ;
        RECT 3.71 1.2 3.8 1.48 ;
        RECT 1.82 1.085 1.91 1.48 ;
        RECT 0.07 0.855 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5 0.08 ;
        RECT 4.755 -0.08 4.845 0.375 ;
        RECT 4.24 -0.08 4.33 0.36 ;
        RECT 3.7 -0.08 3.79 0.36 ;
        RECT 1.805 -0.08 1.895 0.33 ;
        RECT 0.045 -0.08 0.185 0.32 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.555 0.545 0.78 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.425 0.175 0.65 ;
      LAYER MET2 ;
        RECT 0.05 0.23 0.15 0.76 ;
      LAYER VIA1 ;
        RECT 0.055 0.455 0.145 0.545 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.658 0.53 3.02 0.62 ;
        RECT 2.553 0.511 2.696 0.534 ;
        RECT 1.555 0.481 2.658 0.515 ;
        RECT 2.637 0.53 3.02 0.61 ;
        RECT 1.555 0.448 2.637 0.515 ;
        RECT 2.591 0.53 3.02 0.576 ;
        RECT 1.555 0.425 2.591 0.515 ;
        RECT 2.02 0.425 2.28 0.56 ;
      LAYER MET2 ;
        RECT 2.05 0.23 2.15 0.76 ;
      LAYER VIA1 ;
        RECT 2.055 0.455 2.145 0.545 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.975 0.225 4.145 0.375 ;
        RECT 3.975 0.225 4.065 0.92 ;
      LAYER MET2 ;
        RECT 4.05 0.18 4.15 0.56 ;
      LAYER VIA1 ;
        RECT 4.055 0.255 4.145 0.345 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.505 0.25 4.595 0.92 ;
        RECT 4.42 0.25 4.595 0.345 ;
      LAYER MET2 ;
        RECT 4.45 0.18 4.55 0.56 ;
      LAYER VIA1 ;
        RECT 4.455 0.255 4.545 0.345 ;
    END
  END S
  OBS
    LAYER MET1 ;
      RECT 3.795 1.01 4.245 1.1 ;
      RECT 4.155 0.515 4.245 1.1 ;
      RECT 3.795 0.54 3.885 1.1 ;
      RECT 2.485 0.82 2.625 0.91 ;
      RECT 2.485 0.82 2.627 0.909 ;
      RECT 2.485 0.82 2.665 0.889 ;
      RECT 3.16 0.35 3.25 0.87 ;
      RECT 2.587 0.801 3.25 0.87 ;
      RECT 2.627 0.78 3.25 0.87 ;
      RECT 2.625 0.781 3.25 0.87 ;
      RECT 4.155 0.515 4.395 0.655 ;
      RECT 3.16 0.54 3.885 0.63 ;
      RECT 2.734 0.35 3.25 0.44 ;
      RECT 2.713 0.301 2.734 0.43 ;
      RECT 2.667 0.268 2.713 0.396 ;
      RECT 2.629 0.331 2.772 0.354 ;
      RECT 2.485 0.245 2.667 0.335 ;
      RECT 2 1.14 3.61 1.23 ;
      RECT 2 0.905 2.09 1.23 ;
      RECT 0.635 1.035 1.73 1.125 ;
      RECT 1.64 0.905 1.73 1.125 ;
      RECT 0.635 0.395 0.725 1.125 ;
      RECT 1.64 0.905 2.09 0.995 ;
      RECT 0.505 0.895 0.725 0.985 ;
      RECT 0.635 0.395 1.315 0.485 ;
      RECT 1.175 0.36 1.315 0.485 ;
      RECT 0.62 0.336 0.635 0.465 ;
      RECT 0.576 0.392 0.686 0.435 ;
      RECT 0.576 0.367 0.681 0.435 ;
      RECT 0.53 0.19 0.62 0.39 ;
      RECT 3.43 0.17 3.52 0.36 ;
      RECT 2.815 0.17 3.52 0.26 ;
      RECT 2.81 0.96 3.52 1.05 ;
      RECT 3.43 0.85 3.52 1.05 ;
      RECT 1.615 0.65 2.374 0.74 ;
      RECT 1.59 0.65 2.376 0.728 ;
      RECT 1.59 0.65 2.414 0.719 ;
      RECT 0.84 0.625 1.628 0.715 ;
      RECT 2.376 0.61 2.52 0.7 ;
      RECT 2.336 0.631 2.52 0.7 ;
      RECT 2.374 0.611 2.376 0.739 ;
      RECT 0.84 0.637 1.653 0.715 ;
      RECT 0.84 0.575 0.93 0.715 ;
      RECT 0.755 0.17 0.895 0.305 ;
      RECT 0.755 0.17 1.565 0.26 ;
      RECT 0.88 0.855 1.55 0.945 ;
      RECT 1.46 0.805 1.55 0.945 ;
  END
END ADDFX2H7R

MACRO ADDHX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDHX1H7R 0 0 ;
  SIZE 4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4 1.48 ;
        RECT 3.475 1.2 3.615 1.48 ;
        RECT 1.645 1.225 1.785 1.48 ;
        RECT 0.845 1.195 0.935 1.48 ;
        RECT 0.32 1.05 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4 0.08 ;
        RECT 3.43 -0.08 3.57 0.175 ;
        RECT 1.355 -0.08 1.445 0.33 ;
        RECT 0.36 -0.08 0.5 0.21 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.098 1.14 1.38 1.23 ;
        RECT 0.991 1.121 1.136 1.146 ;
        RECT 0.991 1.094 1.098 1.146 ;
        RECT 1.083 1.14 1.38 1.223 ;
        RECT 0.945 1.064 1.083 1.1 ;
        RECT 1.037 1.14 1.38 1.192 ;
        RECT 0.945 1.018 1.037 1.1 ;
        RECT 0.901 0.972 0.991 1.055 ;
        RECT 0.855 0.795 0.945 1.01 ;
        RECT 0.705 0.795 0.945 0.885 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.375 0.73 2.515 0.82 ;
        RECT 2.375 0.387 2.465 0.82 ;
        RECT 2.321 0.342 2.421 0.415 ;
        RECT 2.275 0.314 2.375 0.37 ;
        RECT 2.365 0.387 2.465 0.442 ;
        RECT 2.275 0.17 2.365 0.37 ;
        RECT 1.535 0.17 2.365 0.26 ;
        RECT 1.425 0.455 1.625 0.62 ;
        RECT 1.535 0.17 1.625 0.62 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.295 0.16 0.985 ;
      LAYER MET2 ;
        RECT 0.05 0.625 0.15 1.16 ;
      LAYER VIA1 ;
        RECT 0.055 0.855 0.145 0.945 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.76 0.87 3.91 0.96 ;
        RECT 3.82 0.255 3.91 0.96 ;
        RECT 3.625 0.255 3.91 0.345 ;
      LAYER MET2 ;
        RECT 3.65 0.18 3.75 0.56 ;
      LAYER VIA1 ;
        RECT 3.655 0.255 3.745 0.345 ;
    END
  END S
  OBS
    LAYER MET1 ;
      RECT 2.375 0.96 3.045 1.05 ;
      RECT 2.955 0.715 3.045 1.05 ;
      RECT 2.765 0.715 3.045 0.805 ;
      RECT 3.64 0.604 3.73 0.77 ;
      RECT 2.765 0.17 2.855 0.805 ;
      RECT 3.596 0.514 3.64 0.642 ;
      RECT 3.596 0.559 3.686 0.642 ;
      RECT 3.55 0.469 3.596 0.597 ;
      RECT 3.504 0.423 3.55 0.551 ;
      RECT 3.458 0.377 3.504 0.505 ;
      RECT 3.412 0.331 3.458 0.459 ;
      RECT 3.366 0.285 3.412 0.413 ;
      RECT 3.32 0.239 3.366 0.367 ;
      RECT 3.274 0.193 3.32 0.321 ;
      RECT 2.54 0.215 2.855 0.305 ;
      RECT 3.236 0.239 3.366 0.279 ;
      RECT 2.765 0.17 3.274 0.26 ;
      RECT 2.195 1.14 3.314 1.23 ;
      RECT 2.195 1.14 3.36 1.207 ;
      RECT 3.276 1.121 3.406 1.161 ;
      RECT 2.195 0.53 2.285 1.23 ;
      RECT 1.755 1.045 2.285 1.135 ;
      RECT 3.314 1.079 3.41 1.136 ;
      RECT 3.36 1.033 3.456 1.111 ;
      RECT 3.406 1.008 3.41 1.136 ;
      RECT 3.41 0.695 3.5 1.066 ;
      RECT 1.755 0.91 1.845 1.135 ;
      RECT 1.38 0.91 1.845 1 ;
      RECT 1.865 0.53 2.285 0.62 ;
      RECT 1.865 0.35 1.955 0.62 ;
      RECT 1.815 0.35 1.955 0.44 ;
      RECT 3.205 0.49 3.295 0.99 ;
      RECT 3.03 0.49 3.295 0.58 ;
      RECT 3.03 0.35 3.17 0.58 ;
      RECT 1.11 0.71 1.2 0.985 ;
      RECT 2.015 0.71 2.105 0.85 ;
      RECT 1.11 0.71 2.105 0.8 ;
      RECT 1.175 0.3 1.265 0.8 ;
      RECT 1.065 0.3 1.265 0.39 ;
      RECT 0.555 0.995 0.695 1.085 ;
      RECT 0.524 0.921 0.555 1.05 ;
      RECT 0.478 0.883 0.524 1.011 ;
      RECT 0.478 0.989 0.613 1.011 ;
      RECT 0.478 0.96 0.601 1.011 ;
      RECT 0.432 0.837 0.478 0.965 ;
      RECT 0.386 0.791 0.432 0.919 ;
      RECT 0.34 0.745 0.386 0.873 ;
      RECT 0.296 0.3 0.34 0.828 ;
      RECT 0.25 0.3 0.34 0.783 ;
      RECT 0.25 0.3 0.975 0.39 ;
      RECT 0.475 0.53 1.085 0.62 ;
  END
END ADDHX1H7R

MACRO ADDHX1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDHX1P4H7R 0 0 ;
  SIZE 4.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.2 1.48 ;
        RECT 3.57 1.195 3.71 1.48 ;
        RECT 1.785 1.095 1.925 1.48 ;
        RECT 0.96 1.2 1.05 1.48 ;
        RECT 0.43 1.09 0.52 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.2 0.08 ;
        RECT 3.525 -0.08 3.665 0.175 ;
        RECT 1.515 -0.08 1.605 0.33 ;
        RECT 0.455 -0.08 0.595 0.205 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.208 1.14 1.535 1.23 ;
        RECT 1.113 1.121 1.246 1.158 ;
        RECT 1.113 1.1 1.208 1.158 ;
        RECT 1.205 1.14 1.535 1.229 ;
        RECT 1.067 1.076 1.205 1.112 ;
        RECT 1.159 1.14 1.535 1.204 ;
        RECT 1.067 1.03 1.159 1.112 ;
        RECT 1.021 0.984 1.113 1.066 ;
        RECT 0.975 0.938 1.067 1.02 ;
        RECT 0.931 0.892 1.021 0.975 ;
        RECT 0.885 0.655 0.975 0.93 ;
        RECT 0.825 0.655 0.975 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.54 0.419 2.63 0.845 ;
        RECT 2.501 0.377 2.591 0.458 ;
        RECT 2.455 0.17 2.545 0.415 ;
        RECT 1.715 0.17 2.545 0.26 ;
        RECT 1.515 0.53 1.805 0.62 ;
        RECT 1.715 0.17 1.805 0.62 ;
      LAYER MET2 ;
        RECT 2.45 0.18 2.55 0.56 ;
      LAYER VIA1 ;
        RECT 2.455 0.255 2.545 0.345 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.835 0.255 0.975 ;
        RECT 0.055 0.825 0.235 0.975 ;
        RECT 0.145 0.31 0.235 0.975 ;
      LAYER MET2 ;
        RECT 0.05 0.625 0.15 1.16 ;
      LAYER VIA1 ;
        RECT 0.055 0.855 0.145 0.945 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.825 0.855 3.98 0.945 ;
        RECT 3.89 0.34 3.98 0.945 ;
        RECT 3.81 0.34 3.98 0.43 ;
      LAYER MET2 ;
        RECT 3.85 0.63 3.95 1.16 ;
      LAYER VIA1 ;
        RECT 3.855 0.855 3.945 0.945 ;
    END
  END S
  OBS
    LAYER MET1 ;
      RECT 2.515 0.96 3.14 1.05 ;
      RECT 3.05 0.715 3.14 1.05 ;
      RECT 2.905 0.715 3.14 0.805 ;
      RECT 2.905 0.17 2.995 0.805 ;
      RECT 3.71 0.52 3.8 0.685 ;
      RECT 3.701 0.486 3.71 0.61 ;
      RECT 3.665 0.464 3.701 0.592 ;
      RECT 3.619 0.423 3.665 0.551 ;
      RECT 3.619 0.505 3.739 0.551 ;
      RECT 3.573 0.377 3.619 0.505 ;
      RECT 3.527 0.331 3.573 0.459 ;
      RECT 3.481 0.285 3.527 0.413 ;
      RECT 3.435 0.239 3.481 0.367 ;
      RECT 2.68 0.27 2.995 0.36 ;
      RECT 3.389 0.193 3.435 0.321 ;
      RECT 3.351 0.239 3.481 0.279 ;
      RECT 2.905 0.17 3.389 0.26 ;
      RECT 2.335 1.14 3.404 1.23 ;
      RECT 2.335 1.14 3.45 1.207 ;
      RECT 3.366 1.121 3.48 1.169 ;
      RECT 2.335 0.49 2.425 1.23 ;
      RECT 3.404 1.079 3.526 1.131 ;
      RECT 3.45 1.041 3.48 1.169 ;
      RECT 3.48 0.61 3.57 1.086 ;
      RECT 2.05 0.995 2.425 1.085 ;
      RECT 1.52 0.915 2.14 1.005 ;
      RECT 2.015 0.49 2.425 0.58 ;
      RECT 2.015 0.35 2.105 0.58 ;
      RECT 1.965 0.35 2.105 0.44 ;
      RECT 3.3 0.49 3.39 0.97 ;
      RECT 3.17 0.35 3.31 0.58 ;
      RECT 1.225 0.735 1.315 0.985 ;
      RECT 1.225 0.735 2.245 0.825 ;
      RECT 2.155 0.67 2.245 0.825 ;
      RECT 1.335 0.295 1.425 0.825 ;
      RECT 1.175 0.295 1.425 0.385 ;
      RECT 1.155 0.475 1.245 0.645 ;
      RECT 0.595 0.475 0.685 0.645 ;
      RECT 0.595 0.475 1.245 0.565 ;
      RECT 0.651 0.995 0.81 1.085 ;
      RECT 0.645 0.954 0.651 1.082 ;
      RECT 0.599 0.928 0.645 1.056 ;
      RECT 0.553 0.882 0.599 1.01 ;
      RECT 0.553 0.976 0.689 1.01 ;
      RECT 0.507 0.836 0.553 0.964 ;
      RECT 0.461 0.79 0.507 0.918 ;
      RECT 0.415 0.744 0.461 0.872 ;
      RECT 0.371 0.295 0.415 0.827 ;
      RECT 0.325 0.295 0.415 0.782 ;
      RECT 0.325 0.295 1.085 0.385 ;
  END
END ADDHX1P4H7R

MACRO ADDHX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDHX2H7R 0 0 ;
  SIZE 5 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5 1.48 ;
        RECT 4.3 1.07 4.39 1.48 ;
        RECT 2.09 1.09 2.23 1.48 ;
        RECT 1.1 1.105 1.19 1.48 ;
        RECT 0.57 1.155 0.66 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5 0.08 ;
        RECT 4.21 -0.08 4.35 0.305 ;
        RECT 2.44 -0.08 2.58 0.175 ;
        RECT 1.655 -0.08 1.745 0.33 ;
        RECT 0.595 -0.08 0.735 0.19 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.348 1.045 1.725 1.135 ;
        RECT 1.267 1.026 1.386 1.077 ;
        RECT 1.221 0.989 1.348 1.031 ;
        RECT 1.313 1.045 1.725 1.118 ;
        RECT 1.221 0.949 1.313 1.031 ;
        RECT 1.175 0.903 1.267 0.985 ;
        RECT 1.131 0.857 1.221 0.94 ;
        RECT 1.085 0.645 1.175 0.895 ;
        RECT 0.97 0.645 1.175 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.713 0.17 3.29 0.26 ;
        RECT 3.055 0.17 3.145 0.845 ;
        RECT 2.618 0.246 2.751 0.279 ;
        RECT 2.702 0.175 2.713 0.304 ;
        RECT 2.344 0.265 2.702 0.332 ;
        RECT 2.656 0.204 3.29 0.26 ;
        RECT 2.353 0.265 2.656 0.355 ;
        RECT 2.258 0.245 2.393 0.28 ;
        RECT 1.855 0.22 2.353 0.26 ;
        RECT 2.344 0.265 2.656 0.351 ;
        RECT 1.855 0.193 2.344 0.26 ;
        RECT 2.298 0.265 2.702 0.323 ;
        RECT 1.855 0.17 2.298 0.26 ;
        RECT 1.655 0.545 1.945 0.635 ;
        RECT 1.855 0.17 1.945 0.635 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.305 0.345 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.525 0.83 4.745 0.92 ;
        RECT 4.655 0.235 4.745 0.92 ;
        RECT 4.47 0.235 4.745 0.325 ;
      LAYER MET2 ;
        RECT 4.65 0.425 4.75 0.96 ;
      LAYER VIA1 ;
        RECT 4.655 0.655 4.745 0.745 ;
    END
  END S
  OBS
    LAYER MET1 ;
      RECT 3.125 0.96 3.825 1.05 ;
      RECT 3.525 0.17 3.615 1.05 ;
      RECT 4.395 0.415 4.485 0.685 ;
      RECT 4.151 0.415 4.485 0.505 ;
      RECT 4.128 0.365 4.151 0.494 ;
      RECT 4.082 0.331 4.128 0.459 ;
      RECT 4.082 0.396 4.189 0.459 ;
      RECT 4.036 0.285 4.082 0.413 ;
      RECT 3.99 0.239 4.036 0.367 ;
      RECT 3.944 0.193 3.99 0.321 ;
      RECT 3.906 0.239 4.036 0.279 ;
      RECT 3.525 0.17 3.944 0.26 ;
      RECT 2.87 1.14 4.009 1.23 ;
      RECT 2.87 1.14 4.055 1.207 ;
      RECT 3.971 1.121 4.101 1.161 ;
      RECT 2.87 0.445 2.96 1.23 ;
      RECT 4.009 1.079 4.101 1.161 ;
      RECT 2.335 0.995 2.96 1.085 ;
      RECT 4.055 1.033 4.14 1.119 ;
      RECT 4.101 0.99 4.186 1.076 ;
      RECT 4.14 0.595 4.23 1.031 ;
      RECT 1.825 0.91 2.425 1 ;
      RECT 2.1 0.445 2.96 0.535 ;
      RECT 2.795 0.35 2.885 0.535 ;
      RECT 2.1 0.35 2.19 0.535 ;
      RECT 3.96 0.75 4.05 0.93 ;
      RECT 3.775 0.75 4.05 0.84 ;
      RECT 3.775 0.35 3.865 0.84 ;
      RECT 1.39 0.83 1.565 0.92 ;
      RECT 1.475 0.285 1.565 0.92 ;
      RECT 1.475 0.725 2.78 0.815 ;
      RECT 2.69 0.625 2.78 0.815 ;
      RECT 1.315 0.285 1.565 0.375 ;
      RECT 1.295 0.465 1.385 0.66 ;
      RECT 0.69 0.465 0.78 0.645 ;
      RECT 0.69 0.465 1.385 0.555 ;
      RECT 0.721 0.995 0.95 1.085 ;
      RECT 0.709 0.951 0.721 1.079 ;
      RECT 0.663 0.922 0.709 1.05 ;
      RECT 0.617 0.876 0.663 1.004 ;
      RECT 0.617 0.976 0.759 1.004 ;
      RECT 0.571 0.83 0.617 0.958 ;
      RECT 0.525 0.784 0.571 0.912 ;
      RECT 0.481 0.285 0.525 0.867 ;
      RECT 0.435 0.285 0.525 0.822 ;
      RECT 0.435 0.285 1.225 0.375 ;
  END
END ADDHX2H7R

MACRO AND2X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X0P5H7R 0 0 ;
  SIZE 1.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.2 1.48 ;
        RECT 0.56 1.06 0.7 1.48 ;
        RECT 0.045 0.865 0.185 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.2 0.08 ;
        RECT 0.56 -0.08 0.7 0.245 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.42 0.565 0.55 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.585 0.26 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.85 0.31 0.96 0.98 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.295 0.88 0.76 0.97 ;
      RECT 0.67 0.335 0.76 0.97 ;
      RECT 0.045 0.335 0.76 0.425 ;
  END
END AND2X0P5H7R

MACRO AND2X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X0P7H7R 0 0 ;
  SIZE 1.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.2 1.48 ;
        RECT 0.56 1.045 0.7 1.48 ;
        RECT 0.07 0.865 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.2 0.08 ;
        RECT 0.56 -0.08 0.7 0.245 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.575 0.545 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.85 0.31 0.945 1.005 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.295 0.865 0.76 0.955 ;
      RECT 0.67 0.335 0.76 0.955 ;
      RECT 0.045 0.335 0.76 0.425 ;
  END
END AND2X0P7H7R

MACRO AND2X12H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X12H7R 0 0 ;
  SIZE 4.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.2 1.48 ;
        RECT 4.04 0.83 4.13 1.48 ;
        RECT 3.515 1.02 3.655 1.48 ;
        RECT 3.015 1.02 3.155 1.48 ;
        RECT 2.515 1.02 2.655 1.48 ;
        RECT 2.04 0.98 2.13 1.48 ;
        RECT 1.535 1.095 1.675 1.48 ;
        RECT 0.795 1.095 1.135 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.2 0.08 ;
        RECT 4.04 -0.08 4.13 0.345 ;
        RECT 3.515 -0.08 3.655 0.31 ;
        RECT 3.015 -0.08 3.155 0.31 ;
        RECT 2.515 -0.08 2.655 0.31 ;
        RECT 1.81 -0.08 2.1 0.33 ;
        RECT 1.285 -0.08 1.425 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.2 0.655 1.55 0.745 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.265 0.655 1.005 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.265 0.835 3.945 0.925 ;
        RECT 3.855 0.4 3.945 0.925 ;
        RECT 3.79 0.295 3.88 0.49 ;
        RECT 2.29 0.4 3.945 0.49 ;
        RECT 3.29 0.295 3.38 0.49 ;
        RECT 2.79 0.295 2.88 0.49 ;
        RECT 2.29 0.295 2.38 0.49 ;
      LAYER MET2 ;
        RECT 3.85 0.23 3.95 0.76 ;
      LAYER VIA1 ;
        RECT 3.855 0.455 3.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.81 0.605 1.9 1.035 ;
      RECT 0.07 0.445 0.16 1.035 ;
      RECT 0.07 0.905 1.9 0.995 ;
      RECT 1.81 0.605 3.735 0.695 ;
      RECT 0.07 0.445 0.95 0.535 ;
      RECT 0.81 0.35 0.95 0.535 ;
      RECT 0.295 0.35 0.435 0.535 ;
      RECT 1.09 0.395 1.675 0.485 ;
      RECT 1.09 0.17 1.18 0.485 ;
      RECT 0.045 0.17 0.185 0.325 ;
      RECT 0.545 0.17 0.685 0.305 ;
      RECT 0.045 0.17 1.18 0.26 ;
  END
END AND2X12H7R

MACRO AND2X16H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X16H7R 0 0 ;
  SIZE 4.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.8 1.48 ;
        RECT 4.38 1.07 4.47 1.48 ;
        RECT 3.88 1.07 3.97 1.48 ;
        RECT 3.38 1.07 3.47 1.48 ;
        RECT 2.88 1.07 2.97 1.48 ;
        RECT 2.38 1.055 2.47 1.48 ;
        RECT 1.85 1.095 1.99 1.48 ;
        RECT 1.35 1.095 1.49 1.48 ;
        RECT 0.795 1.095 0.935 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.8 0.08 ;
        RECT 4.355 -0.08 4.495 0.31 ;
        RECT 3.855 -0.08 3.995 0.305 ;
        RECT 3.355 -0.08 3.495 0.305 ;
        RECT 2.855 -0.08 2.995 0.305 ;
        RECT 2.355 -0.08 2.495 0.305 ;
        RECT 1.85 -0.08 1.99 0.305 ;
        RECT 1.35 -0.08 1.49 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.265 0.655 2.015 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.29 0.655 1.03 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.605 0.88 4.745 0.97 ;
        RECT 4.655 0.405 4.745 0.97 ;
        RECT 2.605 0.405 4.745 0.495 ;
        RECT 4.13 0.32 4.22 0.495 ;
      LAYER MET2 ;
        RECT 4.65 0.225 4.75 0.76 ;
      LAYER VIA1 ;
        RECT 4.655 0.455 4.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.125 0.786 2.215 1.035 ;
      RECT 0.07 0.44 0.16 1.035 ;
      RECT 0.07 0.905 2.215 0.995 ;
      RECT 2.171 0.741 2.261 0.824 ;
      RECT 2.215 0.696 2.332 0.749 ;
      RECT 2.261 0.656 2.294 0.785 ;
      RECT 2.294 0.64 4.375 0.73 ;
      RECT 0.07 0.44 0.965 0.53 ;
      RECT 0.875 0.39 0.965 0.53 ;
      RECT 0.295 0.35 0.435 0.53 ;
      RECT 1.14 0.395 2.215 0.485 ;
      RECT 2.125 0.31 2.215 0.485 ;
      RECT 1.625 0.325 1.715 0.485 ;
      RECT 1.14 0.17 1.23 0.485 ;
      RECT 0.045 0.17 0.185 0.325 ;
      RECT 0.545 0.17 0.685 0.305 ;
      RECT 0.045 0.17 1.23 0.26 ;
  END
END AND2X16H7R

MACRO AND2X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X1H7R 0 0 ;
  SIZE 1.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.2 1.48 ;
        RECT 0.59 0.985 0.68 1.48 ;
        RECT 0.085 1.165 0.175 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.2 0.08 ;
        RECT 0.545 -0.08 0.685 0.175 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.37 0.445 0.575 0.595 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.585 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.04 0.24 1.145 0.98 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.325 0.805 0.415 0.945 ;
      RECT 0.325 0.805 0.825 0.895 ;
      RECT 0.735 0.265 0.825 0.895 ;
      RECT 0.05 0.265 0.825 0.355 ;
  END
END AND2X1H7R

MACRO AND2X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X1P4H7R 0 0 ;
  SIZE 1.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.2 1.48 ;
        RECT 0.56 1.025 0.7 1.48 ;
        RECT 0.045 0.87 0.185 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.2 0.08 ;
        RECT 0.52 -0.08 0.66 0.245 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.395 0.595 0.575 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.615 0.23 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.305 0.95 0.975 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.295 0.84 0.76 0.93 ;
      RECT 0.67 0.335 0.76 0.93 ;
      RECT 0.045 0.335 0.76 0.425 ;
  END
END AND2X1P4H7R

MACRO AND2X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X2H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.195 0.91 1.285 1.48 ;
        RECT 0.595 1.095 0.685 1.48 ;
        RECT 0.07 0.92 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.195 -0.08 1.285 0.415 ;
        RECT 0.635 -0.08 0.725 0.21 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.515 0.56 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.945 0.655 1.175 0.745 ;
        RECT 0.945 0.275 1.035 1.025 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.32 0.88 0.41 1.06 ;
      RECT 0.32 0.88 0.85 0.97 ;
      RECT 0.76 0.3 0.85 0.97 ;
      RECT 0.045 0.3 0.85 0.39 ;
  END
END AND2X2H7R

MACRO AND2X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X3H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.195 0.92 1.285 1.48 ;
        RECT 0.595 1.045 0.685 1.48 ;
        RECT 0.07 0.92 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.195 -0.08 1.285 0.365 ;
        RECT 0.635 -0.08 0.725 0.21 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.55 0.56 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.945 0.655 1.175 0.745 ;
        RECT 0.945 0.275 1.035 1.025 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.32 0.865 0.41 1.01 ;
      RECT 0.32 0.865 0.85 0.955 ;
      RECT 0.76 0.325 0.85 0.955 ;
      RECT 0.045 0.325 0.85 0.415 ;
  END
END AND2X3H7R

MACRO AND2X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X4H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 1.855 1.13 1.995 1.48 ;
        RECT 1.36 1.035 1.45 1.48 ;
        RECT 0.34 1.075 0.68 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 1.86 -0.08 1.95 0.36 ;
        RECT 1.36 -0.08 1.45 0.375 ;
        RECT 0.84 -0.08 0.98 0.335 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.725 0.655 1.065 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.625 0.545 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.585 0.95 2.245 1.04 ;
        RECT 2.155 0.285 2.245 1.04 ;
        RECT 1.61 0.455 2.245 0.545 ;
        RECT 2.15 0.285 2.245 0.545 ;
        RECT 1.61 0.3 1.7 0.545 ;
      LAYER MET2 ;
        RECT 1.85 0.225 1.95 0.76 ;
      LAYER VIA1 ;
        RECT 1.855 0.455 1.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.885 1.245 0.975 ;
      RECT 1.155 0.675 1.245 0.975 ;
      RECT 0.07 0.43 0.16 0.975 ;
      RECT 1.155 0.675 2.055 0.765 ;
      RECT 0.07 0.43 0.465 0.52 ;
      RECT 0.325 0.35 0.465 0.52 ;
      RECT 0.59 0.425 1.22 0.515 ;
      RECT 1.13 0.225 1.22 0.515 ;
      RECT 0.59 0.17 0.68 0.515 ;
      RECT 0.045 0.17 0.185 0.34 ;
      RECT 0.045 0.17 0.68 0.26 ;
  END
END AND2X4H7R

MACRO AND2X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X6H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 2.13 0.97 2.22 1.48 ;
        RECT 1.605 1.01 1.745 1.48 ;
        RECT 1.09 1.025 1.23 1.48 ;
        RECT 0.56 1.025 0.7 1.48 ;
        RECT 0.07 0.875 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 2.05 -0.08 2.14 0.345 ;
        RECT 1.525 -0.08 1.665 0.305 ;
        RECT 1.05 -0.08 1.14 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.17 0.655 1.03 0.745 ;
        RECT 0.94 0.605 1.03 0.745 ;
        RECT 0.17 0.535 0.26 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.435 0.455 0.775 0.545 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.855 0.395 1.97 0.975 ;
        RECT 1.8 0.295 1.89 0.485 ;
        RECT 1.38 0.82 1.97 0.91 ;
        RECT 1.3 0.395 1.97 0.485 ;
        RECT 1.38 0.82 1.47 0.96 ;
        RECT 1.3 0.295 1.39 0.485 ;
      LAYER MET2 ;
        RECT 1.85 0.625 1.95 1.16 ;
      LAYER VIA1 ;
        RECT 1.855 0.855 1.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.295 0.845 1.21 0.935 ;
      RECT 1.12 0.42 1.21 0.935 ;
      RECT 1.12 0.595 1.745 0.685 ;
      RECT 0.865 0.42 1.21 0.51 ;
      RECT 0.865 0.225 0.955 0.51 ;
      RECT 0.505 0.225 0.955 0.315 ;
  END
END AND2X6H7R

MACRO AND2X8H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X8H7R 0 0 ;
  SIZE 3 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3 1.48 ;
        RECT 2.56 1.095 2.7 1.48 ;
        RECT 2.06 1.095 2.2 1.48 ;
        RECT 1.56 1.095 1.7 1.48 ;
        RECT 0.81 1.095 0.95 1.48 ;
        RECT 0.085 1.055 0.175 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3 0.08 ;
        RECT 2.56 -0.08 2.7 0.325 ;
        RECT 2.06 -0.08 2.2 0.325 ;
        RECT 1.585 -0.08 1.675 0.345 ;
        RECT 1.085 -0.08 1.175 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.075 0.655 1.415 0.745 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.24 0.655 0.58 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.835 0.31 2.925 1.04 ;
        RECT 1.81 0.91 2.925 1 ;
        RECT 1.835 0.455 2.925 0.545 ;
        RECT 2.335 0.325 2.425 0.545 ;
        RECT 1.835 0.325 1.925 0.545 ;
      LAYER MET2 ;
        RECT 2.65 0.23 2.75 0.76 ;
      LAYER VIA1 ;
        RECT 2.655 0.455 2.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.31 0.905 1.68 0.995 ;
      RECT 1.59 0.68 1.68 0.995 ;
      RECT 0.675 0.35 0.765 0.995 ;
      RECT 1.59 0.68 2.725 0.77 ;
      RECT 0.085 0.41 0.765 0.5 ;
      RECT 0.56 0.35 0.765 0.5 ;
      RECT 0.085 0.205 0.175 0.5 ;
      RECT 0.905 0.435 1.425 0.525 ;
      RECT 1.335 0.285 1.425 0.525 ;
      RECT 0.905 0.17 0.995 0.525 ;
      RECT 0.31 0.17 0.45 0.32 ;
      RECT 0.31 0.17 0.995 0.26 ;
  END
END AND2X8H7R

MACRO AND3X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X0P5H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.84 1.08 0.98 1.48 ;
        RECT 0.31 1.08 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.805 -0.08 0.945 0.335 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.425 0.82 0.625 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.225 0.565 0.625 ;
      LAYER MET2 ;
        RECT 0.45 0.18 0.55 0.56 ;
      LAYER VIA1 ;
        RECT 0.455 0.255 0.545 0.345 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.245 0.425 0.345 0.695 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.105 0.9 1.29 0.99 ;
        RECT 1.2 0.225 1.29 0.99 ;
        RECT 1.055 0.225 1.29 0.375 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.56 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.9 1.01 0.99 ;
      RECT 0.92 0.525 1.01 0.99 ;
      RECT 0.045 0.255 0.135 0.99 ;
      RECT 0.92 0.525 1.11 0.615 ;
      RECT 0.045 0.255 0.185 0.345 ;
  END
END AND3X0P5H7R

MACRO AND3X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X0P7H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.855 1.045 0.995 1.48 ;
        RECT 0.325 1.045 0.465 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.85 -0.08 0.94 0.41 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.595 0.805 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.41 0.555 0.68 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.55 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.15 0.225 1.24 1.145 ;
        RECT 1.055 0.225 1.24 0.375 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.56 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.59 0.865 0.73 1.135 ;
      RECT 0.045 0.865 0.2 1.135 ;
      RECT 0.045 0.865 1.06 0.955 ;
      RECT 0.97 0.63 1.06 0.955 ;
      RECT 0.045 0.31 0.135 1.135 ;
      RECT 0.045 0.31 0.2 0.4 ;
  END
END AND3X0P7H7R

MACRO AND3X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X1H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.85 1.025 0.995 1.48 ;
        RECT 0.32 1.025 0.465 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.825 -0.08 0.965 0.34 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.425 0.785 0.635 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.465 0.225 0.555 0.635 ;
        RECT 0.455 0.225 0.555 0.395 ;
      LAYER MET2 ;
        RECT 0.45 0.18 0.55 0.56 ;
      LAYER VIA1 ;
        RECT 0.455 0.255 0.545 0.345 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.565 0.375 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.15 0.225 1.24 1.055 ;
        RECT 1.06 0.225 1.24 0.395 ;
      LAYER MET2 ;
        RECT 1.055 0.18 1.155 0.56 ;
      LAYER VIA1 ;
        RECT 1.06 0.255 1.15 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.59 0.835 0.73 1.1 ;
      RECT 0.045 0.835 0.2 1.1 ;
      RECT 0.045 0.835 1.06 0.925 ;
      RECT 0.97 0.585 1.06 0.925 ;
      RECT 0.045 0.295 0.135 1.1 ;
      RECT 0.045 0.295 0.2 0.385 ;
  END
END AND3X1H7R

MACRO AND3X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X1P4H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.85 1.045 0.995 1.48 ;
        RECT 0.32 1.045 0.465 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.85 -0.08 0.94 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.575 0.79 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.385 0.555 0.655 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.235 0.55 0.355 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.15 0.225 1.24 1.16 ;
        RECT 1.055 0.225 1.24 0.375 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.56 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.59 0.865 0.73 1.16 ;
      RECT 0.055 0.865 0.2 1.135 ;
      RECT 0.055 0.865 1.06 0.955 ;
      RECT 0.97 0.615 1.06 0.955 ;
      RECT 0.055 0.325 0.145 1.135 ;
      RECT 0.055 0.325 0.2 0.415 ;
  END
END AND3X1P4H7R

MACRO AND3X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X2H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.395 0.945 1.485 1.48 ;
        RECT 0.865 1.11 0.955 1.48 ;
        RECT 0.335 1.11 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.41 -0.08 1.5 0.415 ;
        RECT 0.84 -0.08 0.93 0.415 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.625 0.835 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.4 0.565 0.625 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.565 0.35 0.835 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.105 0.985 1.305 1.075 ;
        RECT 1.215 0.485 1.305 1.075 ;
        RECT 1.055 0.485 1.305 0.575 ;
        RECT 1.055 0.27 1.185 0.575 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.93 1.015 1.02 ;
      RECT 0.925 0.7 1.015 1.02 ;
      RECT 0.045 0.265 0.16 1.02 ;
      RECT 0.925 0.7 1.11 0.79 ;
  END
END AND3X2H7R

MACRO AND3X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X3H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.395 1.035 1.485 1.48 ;
        RECT 0.865 1.105 0.955 1.48 ;
        RECT 0.31 1.105 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.41 -0.08 1.5 0.345 ;
        RECT 0.84 -0.08 0.93 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.625 0.835 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.4 0.565 0.625 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.565 0.35 0.835 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.105 0.93 1.305 1.02 ;
        RECT 1.215 0.485 1.305 1.02 ;
        RECT 1.055 0.485 1.305 0.575 ;
        RECT 1.055 0.27 1.185 0.575 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.925 1.015 1.015 ;
      RECT 0.925 0.7 1.015 1.015 ;
      RECT 0.045 0.205 0.16 1.015 ;
      RECT 0.925 0.7 1.11 0.79 ;
  END
END AND3X3H7R

MACRO AND3X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X4H7R 0 0 ;
  SIZE 3 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3 1.48 ;
        RECT 2.76 1.055 2.85 1.48 ;
        RECT 2.235 1.095 2.375 1.48 ;
        RECT 1.735 1.095 1.875 1.48 ;
        RECT 1.235 1.095 1.375 1.48 ;
        RECT 0.56 1.095 0.7 1.48 ;
        RECT 0.085 1.065 0.175 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3 0.08 ;
        RECT 2.76 -0.08 2.85 0.365 ;
        RECT 2.26 -0.08 2.35 0.35 ;
        RECT 1.76 -0.08 1.85 0.35 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.735 1.725 0.825 ;
        RECT 0.055 0.625 0.145 0.825 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.36 0.35 1.45 0.575 ;
        RECT 0.891 0.35 1.45 0.44 ;
        RECT 0.796 0.331 0.929 0.364 ;
        RECT 0.425 0.306 0.891 0.345 ;
        RECT 0.88 0.35 1.45 0.435 ;
        RECT 0.425 0.278 0.88 0.345 ;
        RECT 0.834 0.35 1.45 0.406 ;
        RECT 0.425 0.255 0.834 0.345 ;
        RECT 0.425 0.255 0.515 0.575 ;
      LAYER MET2 ;
        RECT 0.45 0.18 0.55 0.56 ;
      LAYER VIA1 ;
        RECT 0.455 0.255 0.545 0.345 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.53 1.08 0.62 ;
        RECT 0.625 0.455 0.775 0.62 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.51 0.24 2.6 1.14 ;
        RECT 2.01 0.915 2.6 1.005 ;
        RECT 2.01 0.455 2.6 0.545 ;
        RECT 2.01 0.915 2.1 1.14 ;
        RECT 2.01 0.24 2.1 0.545 ;
      LAYER MET2 ;
        RECT 2.45 0.225 2.55 0.76 ;
      LAYER VIA1 ;
        RECT 2.455 0.455 2.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.51 0.915 1.6 1.195 ;
      RECT 0.92 0.915 1.01 1.195 ;
      RECT 0.335 0.915 0.425 1.195 ;
      RECT 0.335 0.915 1.905 1.005 ;
      RECT 1.815 0.555 1.905 1.005 ;
      RECT 1.815 0.735 2.305 0.825 ;
      RECT 1.54 0.555 1.905 0.645 ;
      RECT 1.54 0.17 1.63 0.645 ;
      RECT 0.97 0.17 1.63 0.26 ;
  END
END AND3X4H7R

MACRO AND3X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X6H7R 0 0 ;
  SIZE 3 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3 1.48 ;
        RECT 2.76 1.055 2.85 1.48 ;
        RECT 2.235 1.095 2.375 1.48 ;
        RECT 1.735 1.095 1.875 1.48 ;
        RECT 1.235 1.095 1.375 1.48 ;
        RECT 0.56 1.095 0.7 1.48 ;
        RECT 0.085 1.055 0.175 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3 0.08 ;
        RECT 2.76 -0.08 2.85 0.365 ;
        RECT 2.26 -0.08 2.35 0.35 ;
        RECT 1.76 -0.08 1.85 0.35 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.71 1.725 0.8 ;
        RECT 0.055 0.625 0.17 0.8 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.36 0.35 1.45 0.575 ;
        RECT 0.891 0.35 1.45 0.44 ;
        RECT 0.796 0.331 0.929 0.364 ;
        RECT 0.425 0.306 0.891 0.345 ;
        RECT 0.88 0.35 1.45 0.435 ;
        RECT 0.425 0.278 0.88 0.345 ;
        RECT 0.834 0.35 1.45 0.406 ;
        RECT 0.425 0.255 0.834 0.345 ;
        RECT 0.425 0.255 0.515 0.575 ;
      LAYER MET2 ;
        RECT 0.45 0.18 0.55 0.56 ;
      LAYER VIA1 ;
        RECT 0.455 0.255 0.545 0.345 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.53 1.08 0.62 ;
        RECT 0.625 0.455 0.775 0.62 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.51 0.315 2.6 1.045 ;
        RECT 2.01 0.905 2.6 0.995 ;
        RECT 2.01 0.455 2.6 0.545 ;
        RECT 2.01 0.905 2.1 1.045 ;
        RECT 2.01 0.315 2.1 0.545 ;
      LAYER MET2 ;
        RECT 2.45 0.225 2.55 0.76 ;
      LAYER VIA1 ;
        RECT 2.455 0.455 2.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.51 0.915 1.6 1.14 ;
      RECT 0.92 0.915 1.01 1.14 ;
      RECT 0.335 0.915 0.425 1.14 ;
      RECT 0.335 0.915 1.905 1.005 ;
      RECT 1.815 0.485 1.905 1.005 ;
      RECT 1.815 0.67 2.305 0.76 ;
      RECT 1.54 0.485 1.905 0.575 ;
      RECT 1.54 0.17 1.63 0.575 ;
      RECT 0.97 0.17 1.63 0.26 ;
  END
END AND3X6H7R

MACRO AND3X8H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X8H7R 0 0 ;
  SIZE 3.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.2 1.48 ;
        RECT 2.65 1.075 2.79 1.48 ;
        RECT 2.15 1.075 2.29 1.48 ;
        RECT 1.635 1.215 1.775 1.48 ;
        RECT 1.105 1.215 1.245 1.48 ;
        RECT 0.575 1.215 0.715 1.48 ;
        RECT 0.085 1.035 0.175 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.2 0.08 ;
        RECT 2.675 -0.08 2.765 0.33 ;
        RECT 2.175 -0.08 2.265 0.33 ;
        RECT 1.675 -0.08 1.765 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.185 0.855 1.585 0.945 ;
        RECT 1.495 0.705 1.585 0.945 ;
        RECT 0.185 0.705 0.275 0.945 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.245 0.455 1.335 0.75 ;
        RECT 0.445 0.455 1.335 0.545 ;
        RECT 0.445 0.455 0.535 0.635 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.74 0.655 1.08 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.925 0.295 3.015 1.02 ;
        RECT 1.925 0.895 3.015 0.985 ;
        RECT 1.925 0.455 3.015 0.545 ;
        RECT 2.425 0.31 2.515 0.545 ;
        RECT 1.925 0.895 2.015 1.035 ;
        RECT 1.925 0.31 2.015 0.545 ;
      LAYER MET2 ;
        RECT 2.85 0.23 2.95 0.76 ;
      LAYER VIA1 ;
        RECT 2.855 0.455 2.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.31 1.035 1.765 1.125 ;
      RECT 1.675 0.52 1.765 1.125 ;
      RECT 1.675 0.635 2.645 0.725 ;
      RECT 1.425 0.52 1.765 0.61 ;
      RECT 1.425 0.275 1.515 0.61 ;
      RECT 0.84 0.275 1.515 0.365 ;
  END
END AND3X8H7R

MACRO AND4X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X0P5H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.1 1.055 1.19 1.48 ;
        RECT 0.56 1.08 0.7 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.1 -0.08 1.19 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.95 0.425 1.175 0.545 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.595 0.805 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.385 0.56 0.61 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.55 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.325 1.08 1.545 1.17 ;
        RECT 1.455 0.23 1.545 1.17 ;
        RECT 1.325 0.23 1.545 0.32 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.825 0.865 0.965 1.17 ;
      RECT 0.295 0.865 0.435 1.17 ;
      RECT 0.045 0.865 1.195 0.955 ;
      RECT 1.105 0.64 1.195 0.955 ;
      RECT 0.045 0.23 0.135 0.955 ;
      RECT 1.105 0.64 1.365 0.73 ;
      RECT 0.045 0.23 0.185 0.32 ;
  END
END AND4X0P5H7R

MACRO AND4X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X0P7H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.075 1.06 1.215 1.48 ;
        RECT 0.56 1.06 0.7 1.48 ;
        RECT 0.045 1.06 0.185 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.1 -0.08 1.19 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.95 0.43 1.175 0.55 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.625 0.835 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.385 0.56 0.61 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.55 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.325 1.06 1.545 1.15 ;
        RECT 1.455 0.25 1.545 1.15 ;
        RECT 1.325 0.25 1.545 0.34 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.825 0.865 0.965 1.15 ;
      RECT 0.295 0.865 0.435 1.15 ;
      RECT 0.045 0.865 1.125 0.955 ;
      RECT 1.035 0.64 1.125 0.955 ;
      RECT 0.045 0.23 0.135 0.955 ;
      RECT 1.035 0.64 1.35 0.73 ;
      RECT 0.045 0.23 0.185 0.32 ;
  END
END AND4X0P7H7R

MACRO AND4X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X1H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.1 1.05 1.19 1.48 ;
        RECT 0.56 1.06 0.7 1.48 ;
        RECT 0.045 1.06 0.185 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.1 -0.08 1.19 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.95 0.425 1.175 0.545 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.595 0.805 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.385 0.56 0.61 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.55 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.325 1.06 1.545 1.15 ;
        RECT 1.455 0.29 1.545 1.15 ;
        RECT 1.325 0.29 1.545 0.38 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.825 0.865 0.965 1.15 ;
      RECT 0.295 0.865 0.435 1.15 ;
      RECT 0.045 0.865 1.125 0.955 ;
      RECT 1.035 0.64 1.125 0.955 ;
      RECT 0.045 0.23 0.135 0.955 ;
      RECT 1.035 0.64 1.365 0.73 ;
      RECT 0.045 0.23 0.185 0.32 ;
  END
END AND4X1H7R

MACRO AND4X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X1P4H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.105 1.06 1.245 1.48 ;
        RECT 0.56 1.06 0.7 1.48 ;
        RECT 0.045 1.06 0.185 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.1 -0.08 1.19 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.95 0.425 1.175 0.545 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.625 0.835 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.385 0.56 0.61 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.55 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.355 1.06 1.545 1.15 ;
        RECT 1.455 0.325 1.545 1.15 ;
        RECT 1.355 0.325 1.545 0.415 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.825 0.865 0.965 1.15 ;
      RECT 0.295 0.865 0.435 1.15 ;
      RECT 0.045 0.865 1.155 0.955 ;
      RECT 1.065 0.64 1.155 0.955 ;
      RECT 0.045 0.24 0.135 0.955 ;
      RECT 1.065 0.64 1.35 0.73 ;
      RECT 0.045 0.24 0.185 0.33 ;
  END
END AND4X1P4H7R

MACRO AND4X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X2H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.64 1.035 1.73 1.48 ;
        RECT 1.1 1.06 1.24 1.48 ;
        RECT 0.56 1.06 0.7 1.48 ;
        RECT 0.045 1.06 0.185 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.64 -0.08 1.73 0.345 ;
        RECT 1.1 -0.08 1.19 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.425 1.145 0.575 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.625 0.835 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.35 0.565 0.575 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.55 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.35 1.06 1.545 1.15 ;
        RECT 1.455 0.245 1.545 1.15 ;
        RECT 1.35 0.245 1.545 0.335 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.825 0.865 0.965 1.15 ;
      RECT 0.295 0.865 0.435 1.15 ;
      RECT 0.045 0.865 1.155 0.955 ;
      RECT 1.065 0.685 1.155 0.955 ;
      RECT 0.045 0.25 0.135 0.955 ;
      RECT 1.065 0.685 1.365 0.775 ;
      RECT 1.275 0.615 1.365 0.775 ;
      RECT 0.045 0.25 0.185 0.34 ;
  END
END AND4X2H7R

MACRO AND4X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X3H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.64 1.035 1.73 1.48 ;
        RECT 1.075 1.06 1.215 1.48 ;
        RECT 0.555 1.06 0.695 1.48 ;
        RECT 0.045 1.045 0.185 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.64 -0.08 1.73 0.345 ;
        RECT 1.1 -0.08 1.19 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.425 1.145 0.575 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.625 0.835 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.395 0.56 0.62 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.55 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.35 1.06 1.545 1.15 ;
        RECT 1.455 0.32 1.545 1.15 ;
        RECT 1.35 0.32 1.545 0.41 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.825 0.865 0.965 1.15 ;
      RECT 0.295 0.865 0.435 1.15 ;
      RECT 0.045 0.865 1.155 0.955 ;
      RECT 1.065 0.665 1.155 0.955 ;
      RECT 0.045 0.23 0.135 0.955 ;
      RECT 1.065 0.665 1.365 0.755 ;
      RECT 1.275 0.6 1.365 0.755 ;
      RECT 0.045 0.23 0.185 0.32 ;
  END
END AND4X3H7R

MACRO AND4X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X4H7R 0 0 ;
  SIZE 4.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.2 1.48 ;
        RECT 3.885 1.06 4.025 1.48 ;
        RECT 3.355 1.06 3.495 1.48 ;
        RECT 2.8 1.035 2.89 1.48 ;
        RECT 2.53 1.075 2.67 1.48 ;
        RECT 1.955 1.075 2.095 1.48 ;
        RECT 1.165 1.075 1.505 1.48 ;
        RECT 0.575 1.075 0.715 1.48 ;
        RECT 0.085 1.05 0.175 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.2 0.08 ;
        RECT 3.885 -0.08 4.025 0.375 ;
        RECT 3.305 -0.08 3.445 0.375 ;
        RECT 2.81 -0.08 2.9 0.4 ;
        RECT 0.335 -0.08 0.425 0.35 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.21 0.655 0.55 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.74 0.655 1.08 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.56 0.655 1.905 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.155 0.655 2.495 0.745 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.05 0.88 3.945 0.97 ;
        RECT 3.855 0.52 3.945 0.97 ;
        RECT 3.04 0.52 3.945 0.61 ;
        RECT 3.62 0.88 3.76 1.12 ;
        RECT 3.6 0.285 3.74 0.61 ;
        RECT 3.05 0.88 3.19 1.12 ;
        RECT 3.04 0.285 3.18 0.61 ;
      LAYER MET2 ;
        RECT 3.85 0.43 3.95 0.96 ;
      LAYER VIA1 ;
        RECT 3.855 0.655 3.945 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.65 0.895 1.79 1.17 ;
      RECT 0.84 0.895 0.98 1.17 ;
      RECT 2.245 0.895 2.385 1.165 ;
      RECT 0.31 0.895 0.45 1.165 ;
      RECT 0.31 0.895 2.695 0.985 ;
      RECT 2.605 0.445 2.695 0.985 ;
      RECT 2.605 0.7 3.705 0.79 ;
      RECT 2.25 0.445 2.695 0.535 ;
      RECT 2.25 0.355 2.39 0.535 ;
      RECT 2.525 0.175 2.67 0.34 ;
      RECT 1.94 0.175 2.08 0.34 ;
      RECT 1.38 0.175 1.52 0.34 ;
      RECT 1.38 0.175 2.67 0.265 ;
      RECT 0.87 0.435 1.8 0.525 ;
      RECT 1.655 0.355 1.8 0.525 ;
      RECT 0.87 0.35 1.01 0.525 ;
      RECT 0.085 0.44 0.675 0.53 ;
      RECT 0.585 0.17 0.675 0.53 ;
      RECT 0.085 0.225 0.175 0.53 ;
      RECT 1.12 0.17 1.29 0.34 ;
      RECT 0.585 0.17 1.29 0.26 ;
  END
END AND4X4H7R

MACRO AND4X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X6H7R 0 0 ;
  SIZE 4.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.2 1.48 ;
        RECT 3.87 0.965 4.01 1.48 ;
        RECT 3.34 0.965 3.48 1.48 ;
        RECT 2.785 0.92 2.875 1.48 ;
        RECT 2.53 1.06 2.67 1.48 ;
        RECT 1.94 1.06 2.08 1.48 ;
        RECT 1.15 1.06 1.49 1.48 ;
        RECT 0.56 1.06 0.7 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.2 0.08 ;
        RECT 3.87 -0.08 4.01 0.25 ;
        RECT 3.305 -0.08 3.445 0.25 ;
        RECT 2.795 -0.08 2.885 0.365 ;
        RECT 0.32 -0.08 0.41 0.35 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.195 0.655 0.535 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.755 0.655 1.095 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.545 0.655 1.89 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.135 0.655 2.475 0.745 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.06 0.775 3.945 0.865 ;
        RECT 3.855 0.34 3.945 0.865 ;
        RECT 3.02 0.34 3.945 0.43 ;
        RECT 3.63 0.775 3.72 0.915 ;
        RECT 3.06 0.775 3.15 0.915 ;
      LAYER MET2 ;
        RECT 3.85 0.43 3.95 0.96 ;
      LAYER VIA1 ;
        RECT 3.855 0.655 3.945 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.23 0.88 2.37 1.15 ;
      RECT 1.635 0.88 1.775 1.15 ;
      RECT 0.85 0.88 0.99 1.15 ;
      RECT 0.295 0.88 0.435 1.15 ;
      RECT 0.295 0.88 2.655 0.97 ;
      RECT 2.565 0.445 2.655 0.97 ;
      RECT 2.565 0.57 3.69 0.66 ;
      RECT 2.235 0.445 2.655 0.535 ;
      RECT 2.235 0.36 2.375 0.535 ;
      RECT 2.515 0.175 2.655 0.34 ;
      RECT 1.365 0.175 1.505 0.34 ;
      RECT 1.925 0.175 2.065 0.325 ;
      RECT 1.365 0.175 2.655 0.265 ;
      RECT 0.855 0.435 1.785 0.525 ;
      RECT 1.645 0.355 1.785 0.525 ;
      RECT 0.855 0.35 0.995 0.525 ;
      RECT 0.07 0.44 0.66 0.53 ;
      RECT 0.57 0.17 0.66 0.53 ;
      RECT 0.07 0.225 0.16 0.53 ;
      RECT 1.135 0.17 1.275 0.34 ;
      RECT 0.57 0.17 1.275 0.26 ;
  END
END AND4X6H7R

MACRO ANT2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ANT2H7R 0 0 ;
  SIZE 0.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.4 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.4 0.08 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.065 0.425 0.35 0.575 ;
        RECT 0.065 0.28 0.22 1.12 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END A
END ANT2H7R

MACRO ANT4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ANT4H7R 0 0 ;
  SIZE 0.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.8 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.8 0.08 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.062 0.279 0.614 1.12 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END A
END ANT4H7R

MACRO AO211X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO211X0P5H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.34 0.88 1.43 1.48 ;
        RECT 0.845 1.11 0.935 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.1 -0.08 1.24 0.175 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.455 1.25 0.575 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.705 0.655 0.975 0.755 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.55 0.57 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.69 0.345 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.615 0.265 1.745 0.98 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.265 0.16 1.045 ;
      RECT 1.425 0.265 1.515 0.59 ;
      RECT 0.6 0.265 0.69 0.405 ;
      RECT 0.07 0.265 1.515 0.355 ;
      RECT 0.555 0.93 1.225 1.02 ;
  END
END AO211X0P5H7R

MACRO AO211X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO211X0P7H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.34 0.912 1.43 1.48 ;
        RECT 0.845 1.11 0.935 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.1 -0.08 1.24 0.175 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.455 1.25 0.575 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.705 0.655 0.975 0.755 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.55 0.57 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.69 0.345 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.615 0.265 1.745 0.98 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.265 0.16 1.045 ;
      RECT 1.425 0.265 1.515 0.59 ;
      RECT 0.07 0.265 1.515 0.365 ;
      RECT 0.555 0.93 1.225 1.02 ;
  END
END AO211X0P7H7R

MACRO AO211X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO211X1H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.34 0.96 1.43 1.48 ;
        RECT 0.845 1.11 0.935 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.1 -0.08 1.24 0.185 ;
        RECT 0.31 -0.08 0.45 0.185 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.455 1.25 0.575 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.705 0.655 0.975 0.755 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.55 0.57 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.69 0.345 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.615 0.265 1.745 0.98 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.265 0.16 1.045 ;
      RECT 1.425 0.275 1.515 0.59 ;
      RECT 0.07 0.275 1.515 0.365 ;
      RECT 0.555 0.93 1.225 1.02 ;
  END
END AO211X1H7R

MACRO AO211X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO211X1P4H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.34 1.004 1.43 1.48 ;
        RECT 0.845 1.11 0.935 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.1 -0.08 1.24 0.185 ;
        RECT 0.31 -0.08 0.45 0.185 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.455 1.25 0.575 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.705 0.655 0.975 0.755 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.55 0.57 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.69 0.345 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.615 0.301 1.745 0.98 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.265 0.16 1.045 ;
      RECT 1.425 0.275 1.515 0.626 ;
      RECT 0.07 0.275 1.515 0.365 ;
      RECT 0.555 0.93 1.225 1.02 ;
  END
END AO211X1P4H7R

MACRO AO211X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO211X2H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.84 0.97 1.93 1.48 ;
        RECT 1.34 0.97 1.43 1.48 ;
        RECT 0.335 1.135 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.84 -0.08 1.93 0.39 ;
        RECT 1.32 -0.08 1.41 0.375 ;
        RECT 0.56 -0.08 0.7 0.185 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.35 0.455 0.575 0.575 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.625 0.775 0.85 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.93 0.455 1.02 0.65 ;
        RECT 0.825 0.455 1.02 0.545 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.59 0.225 1.745 0.375 ;
        RECT 1.59 0.225 1.68 1.055 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.56 ;
      LAYER VIA1 ;
        RECT 1.655 0.255 1.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.11 0.275 1.2 1.07 ;
      RECT 1.11 0.575 1.48 0.665 ;
      RECT 0.045 0.275 1.2 0.365 ;
      RECT 0.045 0.955 0.715 1.045 ;
  END
END AO211X2H7R

MACRO AO211X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO211X3H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.84 1.055 1.93 1.48 ;
        RECT 1.34 1.055 1.43 1.48 ;
        RECT 0.335 1.135 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.84 -0.08 1.93 0.345 ;
        RECT 1.34 -0.08 1.43 0.33 ;
        RECT 0.56 -0.08 0.7 0.185 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.42 0.455 0.575 0.545 ;
        RECT 0.42 0.455 0.54 0.655 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.625 0.775 0.85 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.93 0.455 1.02 0.65 ;
        RECT 0.825 0.455 1.02 0.545 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.59 0.225 1.745 0.375 ;
        RECT 1.59 0.225 1.68 1.045 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.56 ;
      LAYER VIA1 ;
        RECT 1.655 0.255 1.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.11 0.275 1.2 1.075 ;
      RECT 1.11 0.575 1.48 0.665 ;
      RECT 0.045 0.275 1.2 0.365 ;
      RECT 0.045 0.955 0.715 1.045 ;
  END
END AO211X3H7R

MACRO AO211X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO211X4H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.84 0.855 1.93 1.48 ;
        RECT 1.34 0.855 1.43 1.48 ;
        RECT 0.31 1.075 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.784 -0.08 1.88 0.081 ;
        RECT 1.784 -0.08 1.874 0.345 ;
        RECT 1.279 -0.08 1.369 0.33 ;
        RECT 0.56 -0.08 0.7 0.185 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.455 0.575 0.545 ;
        RECT 0.425 0.455 0.53 0.705 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.655 0.825 0.79 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.93 0.455 1.02 0.705 ;
        RECT 0.825 0.455 1.02 0.545 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.59 0.655 1.775 0.745 ;
        RECT 1.59 0.395 1.68 1.15 ;
        RECT 1.509 0.395 1.68 0.485 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.11 0.356 1.2 1.015 ;
      RECT 1.11 0.65 1.48 0.74 ;
      RECT 1.097 0.281 1.11 0.41 ;
      RECT 1.059 0.356 1.2 0.384 ;
      RECT 0.045 0.275 1.097 0.365 ;
      RECT 0.045 0.311 1.156 0.365 ;
      RECT 0.045 0.895 0.185 1.015 ;
      RECT 0.045 0.895 0.705 0.985 ;
  END
END AO211X4H7R

MACRO AO211X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO211X6H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 2.147 1.055 2.237 1.48 ;
        RECT 1.647 0.855 1.737 1.48 ;
        RECT 0.527 1.095 0.667 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 1.907 -0.08 2.047 0.305 ;
        RECT 1.432 -0.08 1.522 0.33 ;
        RECT 0.842 -0.08 0.982 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.702 0.455 0.792 0.705 ;
        RECT 0.625 0.455 0.792 0.545 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.397 0.625 0.577 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.915 0.625 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.615 1.372 0.975 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.397 0.395 2.487 1.165 ;
        RECT 1.897 0.855 2.487 0.945 ;
        RECT 1.657 0.395 2.487 0.485 ;
        RECT 2.182 0.225 2.272 0.485 ;
        RECT 1.897 0.855 1.987 1.195 ;
      LAYER MET2 ;
        RECT 2.25 0.63 2.35 1.16 ;
      LAYER VIA1 ;
        RECT 2.255 0.855 2.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.357 1.08 1.557 1.17 ;
      RECT 1.467 0.435 1.557 1.17 ;
      RECT 1.467 0.63 1.927 0.72 ;
      RECT 1.207 0.435 1.557 0.525 ;
      RECT 1.207 0.275 1.297 0.525 ;
      RECT 0.297 0.275 1.297 0.365 ;
      RECT 0.781 0.88 0.921 1.17 ;
      RECT 0.277 0.88 0.417 1.17 ;
      RECT 0.277 0.88 0.921 0.97 ;
  END
END AO211X6H7R

MACRO AO21X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21X0P5H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.11 0.845 1.2 1.48 ;
        RECT 0.31 1.05 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.87 -0.08 1.01 0.175 ;
        RECT 0.07 -0.08 0.16 0.37 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.595 0.205 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.425 0.545 0.725 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.575 0.79 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.385 0.254 1.475 0.945 ;
        RECT 1.225 0.254 1.475 0.345 ;
      LAYER MET2 ;
        RECT 1.25 0.18 1.35 0.56 ;
      LAYER VIA1 ;
        RECT 1.255 0.255 1.345 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.88 0.265 0.97 0.95 ;
      RECT 0.88 0.575 1.295 0.665 ;
      RECT 0.605 0.265 0.97 0.355 ;
      RECT 0.045 0.87 0.715 0.96 ;
  END
END AO21X0P5H7R

MACRO AO21X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21X0P7H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.11 0.877 1.2 1.48 ;
        RECT 0.31 1.045 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.87 -0.08 1.01 0.175 ;
        RECT 0.07 -0.08 0.16 0.37 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.595 0.205 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.425 0.545 0.725 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.575 0.79 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.385 0.254 1.475 0.945 ;
        RECT 1.225 0.254 1.475 0.345 ;
      LAYER MET2 ;
        RECT 1.25 0.18 1.35 0.56 ;
      LAYER VIA1 ;
        RECT 1.255 0.255 1.345 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.88 0.265 0.97 0.945 ;
      RECT 0.88 0.575 1.295 0.665 ;
      RECT 0.605 0.265 0.97 0.355 ;
      RECT 0.045 0.865 0.715 0.955 ;
  END
END AO21X0P7H7R

MACRO AO21X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21X1H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.125 0.925 1.215 1.48 ;
        RECT 0.31 1.05 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.87 -0.08 1.01 0.175 ;
        RECT 0.07 -0.08 0.16 0.37 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.595 0.205 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.425 0.545 0.725 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.595 0.805 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.385 0.255 1.475 0.975 ;
        RECT 1.225 0.255 1.475 0.346 ;
      LAYER MET2 ;
        RECT 1.25 0.18 1.35 0.56 ;
      LAYER VIA1 ;
        RECT 1.255 0.255 1.345 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.895 0.265 0.985 0.95 ;
      RECT 0.895 0.575 1.295 0.665 ;
      RECT 0.605 0.265 0.985 0.355 ;
      RECT 0.045 0.87 0.715 0.96 ;
  END
END AO21X1H7R

MACRO AO21X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21X1P4H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.11 0.969 1.2 1.48 ;
        RECT 0.31 1.05 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.87 -0.08 1.01 0.175 ;
        RECT 0.07 -0.08 0.16 0.37 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.595 0.205 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.425 0.545 0.725 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.575 0.79 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.385 0.254 1.475 0.945 ;
        RECT 1.225 0.254 1.475 0.345 ;
      LAYER MET2 ;
        RECT 1.25 0.18 1.35 0.56 ;
      LAYER VIA1 ;
        RECT 1.255 0.255 1.345 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.88 0.265 0.97 0.95 ;
      RECT 0.88 0.575 1.295 0.665 ;
      RECT 0.605 0.265 0.97 0.355 ;
      RECT 0.045 0.87 0.715 0.96 ;
  END
END AO21X1P4H7R

MACRO AO21X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21X2H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.625 0.845 1.715 1.48 ;
        RECT 1.125 0.845 1.215 1.48 ;
        RECT 0.31 1.05 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.555 -0.08 1.645 0.37 ;
        RECT 0.87 -0.08 1.01 0.175 ;
        RECT 0.07 -0.08 0.16 0.37 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.595 0.205 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.425 0.545 0.725 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.595 0.805 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.375 0.254 1.465 0.93 ;
        RECT 1.225 0.254 1.465 0.345 ;
      LAYER MET2 ;
        RECT 1.25 0.18 1.35 0.56 ;
      LAYER VIA1 ;
        RECT 1.255 0.255 1.345 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.895 0.265 0.985 0.945 ;
      RECT 0.895 0.575 1.255 0.665 ;
      RECT 0.605 0.265 0.985 0.355 ;
      RECT 0.045 0.87 0.715 0.96 ;
  END
END AO21X2H7R

MACRO AO21X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21X3H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.625 0.94 1.715 1.48 ;
        RECT 1.125 0.94 1.215 1.48 ;
        RECT 0.31 1.045 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.555 -0.08 1.645 0.37 ;
        RECT 0.87 -0.08 1.01 0.175 ;
        RECT 0.07 -0.08 0.16 0.37 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.595 0.205 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.425 0.545 0.725 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.595 0.805 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.375 0.254 1.465 0.93 ;
        RECT 1.225 0.254 1.465 0.345 ;
      LAYER MET2 ;
        RECT 1.25 0.18 1.35 0.56 ;
      LAYER VIA1 ;
        RECT 1.255 0.255 1.345 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.895 0.265 0.985 0.945 ;
      RECT 0.895 0.575 1.255 0.665 ;
      RECT 0.605 0.265 0.985 0.355 ;
      RECT 0.045 0.865 0.715 0.955 ;
  END
END AO21X3H7R

MACRO AO21X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21X4H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.595 1.055 1.685 1.48 ;
        RECT 1.095 1.055 1.185 1.48 ;
        RECT 0.31 1.07 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.51 -0.08 1.6 0.345 ;
        RECT 0.82 -0.08 0.96 0.175 ;
        RECT 0.07 -0.08 0.16 0.35 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.595 0.205 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.425 0.545 0.695 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.575 0.775 0.8 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.225 0.855 1.435 0.95 ;
        RECT 1.345 0.395 1.435 0.95 ;
        RECT 1.135 0.395 1.435 0.485 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.865 0.434 0.955 1.005 ;
      RECT 0.865 0.625 1.205 0.715 ;
      RECT 0.836 0.351 0.865 0.48 ;
      RECT 0.79 0.314 0.836 0.442 ;
      RECT 0.79 0.389 0.911 0.442 ;
      RECT 0.744 0.268 0.79 0.396 ;
      RECT 0.706 0.245 0.744 0.354 ;
      RECT 0.505 0.245 0.744 0.335 ;
      RECT 0.045 0.89 0.715 0.98 ;
  END
END AO21X4H7R

MACRO AO21X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21X6H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 1.907 1.07 1.997 1.48 ;
        RECT 1.407 1.055 1.497 1.48 ;
        RECT 0.588 1.07 0.678 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 1.651 -0.08 1.791 0.305 ;
        RECT 1.126 -0.08 1.216 0.33 ;
        RECT 0.323 -0.08 0.413 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.625 0.476 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.425 0.765 0.705 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.615 1.046 0.795 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.591 0.855 2.272 0.945 ;
        RECT 1.998 0.301 2.088 0.945 ;
        RECT 1.401 0.395 2.088 0.485 ;
        RECT 1.901 0.301 2.088 0.485 ;
      LAYER MET2 ;
        RECT 2.05 0.63 2.15 1.16 ;
      LAYER VIA1 ;
        RECT 2.055 0.855 2.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.136 0.435 1.226 0.965 ;
      RECT 1.136 0.625 1.908 0.715 ;
      RECT 0.876 0.435 1.226 0.525 ;
      RECT 0.876 0.37 0.966 0.525 ;
      RECT 0.298 0.89 0.968 0.98 ;
  END
END AO21X6H7R

MACRO AO21X8H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21X8H7R 0 0 ;
  SIZE 3.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.6 1.48 ;
        RECT 3.075 1.055 3.165 1.48 ;
        RECT 2.575 1.07 2.665 1.48 ;
        RECT 2.075 1.055 2.165 1.48 ;
        RECT 1.04 1.015 1.18 1.48 ;
        RECT 0.31 1.015 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.6 0.08 ;
        RECT 3.075 -0.08 3.165 0.345 ;
        RECT 2.55 -0.08 2.69 0.305 ;
        RECT 2.075 -0.08 2.165 0.345 ;
        RECT 1.57 -0.08 1.71 0.31 ;
        RECT 0.575 -0.08 0.715 0.325 ;
        RECT 0.1 -0.08 0.19 0.35 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.195 0.655 0.535 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.89 0.655 1.23 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.445 0.655 1.785 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.3 0.855 2.945 0.945 ;
        RECT 2.855 0.395 2.945 0.945 ;
        RECT 2.3 0.395 2.945 0.485 ;
      LAYER MET2 ;
        RECT 2.85 0.43 2.95 0.96 ;
      LAYER VIA1 ;
        RECT 2.855 0.655 2.945 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.555 0.865 1.965 0.955 ;
      RECT 1.875 0.335 1.965 0.955 ;
      RECT 1.875 0.625 2.765 0.715 ;
      RECT 1.345 0.4 1.965 0.49 ;
      RECT 1.82 0.335 1.965 0.49 ;
      RECT 1.345 0.17 1.435 0.49 ;
      RECT 0.805 0.17 0.945 0.325 ;
      RECT 0.805 0.17 1.435 0.26 ;
      RECT 1.33 1.045 1.96 1.135 ;
      RECT 1.33 0.835 1.42 1.135 ;
      RECT 0.07 0.835 0.16 0.975 ;
      RECT 0.07 0.835 1.42 0.925 ;
      RECT 0.35 0.415 1.195 0.505 ;
      RECT 1.055 0.35 1.195 0.505 ;
      RECT 0.35 0.325 0.44 0.505 ;
  END
END AO21X8H7R

MACRO AO221X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO221X0P5H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.79 0.82 1.88 1.48 ;
        RECT 0.54 1.215 0.63 1.48 ;
        RECT 0.085 1.215 0.175 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.765 -0.08 1.855 0.35 ;
        RECT 0.64 -0.08 0.78 0.16 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.455 0.585 0.635 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.78 0.625 0.96 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.455 1.295 0.555 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.225 0.655 1.495 0.765 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.04 0.225 2.145 0.92 ;
      LAYER MET2 ;
        RECT 2.05 0.18 2.15 0.56 ;
      LAYER VIA1 ;
        RECT 2.055 0.255 2.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.535 0.87 1.675 0.96 ;
      RECT 1.585 0.25 1.675 0.96 ;
      RECT 1.585 0.57 1.95 0.66 ;
      RECT 0.045 0.25 1.675 0.34 ;
      RECT 0.76 1.045 1.39 1.135 ;
      RECT 1.3 0.9 1.39 1.135 ;
      RECT 0.28 0.865 1.165 0.955 ;
  END
END AO221X0P5H7R

MACRO AO221X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO221X0P7H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.79 0.82 1.88 1.48 ;
        RECT 0.54 1.215 0.63 1.48 ;
        RECT 0.085 1.215 0.175 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.765 -0.08 1.855 0.35 ;
        RECT 0.64 -0.08 0.78 0.16 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.455 0.585 0.635 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.78 0.625 0.96 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.455 1.295 0.555 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.225 0.655 1.495 0.765 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.04 0.225 2.145 0.92 ;
      LAYER MET2 ;
        RECT 2.05 0.18 2.15 0.56 ;
      LAYER VIA1 ;
        RECT 2.055 0.255 2.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.535 0.87 1.675 0.96 ;
      RECT 1.585 0.25 1.675 0.96 ;
      RECT 1.585 0.57 1.95 0.66 ;
      RECT 0.045 0.25 1.675 0.34 ;
      RECT 0.76 1.045 1.39 1.135 ;
      RECT 1.3 0.9 1.39 1.135 ;
      RECT 0.28 0.865 1.165 0.955 ;
  END
END AO221X0P7H7R

MACRO AO221X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO221X1H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.79 0.82 1.88 1.48 ;
        RECT 0.54 1.215 0.63 1.48 ;
        RECT 0.085 1.215 0.175 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.765 -0.08 1.855 0.35 ;
        RECT 0.64 -0.08 0.78 0.16 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.455 0.585 0.635 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.78 0.625 0.96 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.455 1.295 0.555 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.225 0.655 1.495 0.765 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.04 0.225 2.145 0.92 ;
      LAYER MET2 ;
        RECT 2.05 0.18 2.15 0.56 ;
      LAYER VIA1 ;
        RECT 2.055 0.255 2.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.535 0.87 1.675 0.96 ;
      RECT 1.585 0.25 1.675 0.96 ;
      RECT 1.585 0.57 1.95 0.66 ;
      RECT 0.045 0.25 1.675 0.34 ;
      RECT 0.76 1.045 1.39 1.135 ;
      RECT 1.3 0.9 1.39 1.135 ;
      RECT 0.28 0.865 1.165 0.955 ;
  END
END AO221X1H7R

MACRO AO221X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO221X1P4H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.79 0.82 1.88 1.48 ;
        RECT 0.54 1.215 0.63 1.48 ;
        RECT 0.085 1.215 0.175 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.765 -0.08 1.855 0.35 ;
        RECT 0.64 -0.08 0.78 0.16 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.455 0.585 0.635 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.78 0.625 0.96 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.455 1.295 0.555 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.225 0.655 1.495 0.765 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.04 0.225 2.145 0.92 ;
      LAYER MET2 ;
        RECT 2.05 0.18 2.15 0.56 ;
      LAYER VIA1 ;
        RECT 2.055 0.255 2.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.535 0.87 1.675 0.96 ;
      RECT 1.585 0.25 1.675 0.96 ;
      RECT 1.585 0.57 1.95 0.66 ;
      RECT 0.07 0.25 1.675 0.345 ;
      RECT 1.3 0.205 1.39 0.345 ;
      RECT 0.07 0.205 0.16 0.345 ;
      RECT 0.76 1.045 1.39 1.135 ;
      RECT 1.3 0.9 1.39 1.135 ;
      RECT 0.28 0.865 1.165 0.955 ;
  END
END AO221X1P4H7R

MACRO AO221X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO221X2H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 1.09 1.225 1.23 1.48 ;
        RECT 0.6 0.905 0.69 1.48 ;
        RECT 0.07 0.905 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 2.115 -0.08 2.255 0.175 ;
        RECT 1.335 -0.08 1.475 0.175 ;
        RECT 0.59 -0.08 0.73 0.175 ;
        RECT 0.07 -0.08 0.16 0.39 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.705 0.655 0.975 0.755 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.455 1.215 0.565 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.385 0.455 1.595 0.545 ;
        RECT 1.385 0.455 1.565 0.6 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.655 0.625 1.835 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.975 0.615 2.145 0.775 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.32 0.225 0.41 1.045 ;
        RECT 0.255 0.225 0.41 0.375 ;
      LAYER MET2 ;
        RECT 0.25 0.18 0.35 0.56 ;
      LAYER VIA1 ;
        RECT 0.255 0.255 0.345 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.24 0.275 2.33 0.98 ;
      RECT 0.5 0.275 0.59 0.675 ;
      RECT 0.5 0.275 2.33 0.365 ;
      RECT 0.85 1.045 1.725 1.135 ;
      RECT 0.85 0.905 0.94 1.135 ;
      RECT 1.32 0.865 1.99 0.955 ;
  END
END AO221X2H7R

MACRO AO221X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO221X3H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 1.09 1.225 1.23 1.48 ;
        RECT 0.58 0.965 0.67 1.48 ;
        RECT 0.07 0.985 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 2.135 -0.08 2.275 0.175 ;
        RECT 1.335 -0.08 1.475 0.175 ;
        RECT 0.59 -0.08 0.73 0.175 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.705 0.655 0.975 0.755 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.02 0.455 1.245 0.575 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.385 0.65 1.61 0.77 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.745 0.455 1.835 0.63 ;
        RECT 1.62 0.455 1.835 0.545 ;
      LAYER MET2 ;
        RECT 1.65 0.23 1.75 0.76 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.975 0.615 2.145 0.775 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.825 0.41 0.975 ;
        RECT 0.32 0.315 0.41 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.24 0.275 2.33 0.98 ;
      RECT 0.5 0.275 0.59 0.65 ;
      RECT 0.5 0.275 2.33 0.365 ;
      RECT 1.075 0.255 1.215 0.365 ;
      RECT 0.85 1.045 1.725 1.135 ;
      RECT 0.85 0.965 0.94 1.135 ;
      RECT 1.32 0.865 2.01 0.955 ;
  END
END AO221X3H7R

MACRO AO221X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO221X4H7R 0 0 ;
  SIZE 2.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.8 1.48 ;
        RECT 1.335 1.225 1.475 1.48 ;
        RECT 0.845 1.05 0.935 1.48 ;
        RECT 0.315 0.855 0.405 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.8 0.08 ;
        RECT 2.38 -0.08 2.52 0.175 ;
        RECT 1.58 -0.08 1.72 0.175 ;
        RECT 0.835 -0.08 0.975 0.175 ;
        RECT 0.295 -0.08 0.385 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.655 1.19 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.285 0.455 1.375 0.65 ;
        RECT 1.18 0.455 1.375 0.545 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.61 0.655 1.835 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.95 0.655 2.175 0.775 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.32 0.455 2.41 0.68 ;
        RECT 2.225 0.455 2.41 0.545 ;
      LAYER MET2 ;
        RECT 2.25 0.23 2.35 0.76 ;
      LAYER VIA1 ;
        RECT 2.255 0.455 2.345 0.545 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.545 1.025 0.745 1.175 ;
        RECT 0.545 0.37 0.655 1.175 ;
      LAYER MET2 ;
        RECT 0.65 0.84 0.75 1.22 ;
      LAYER VIA1 ;
        RECT 0.655 1.055 0.745 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.47 0.845 2.59 0.985 ;
      RECT 2.5 0.275 2.59 0.985 ;
      RECT 0.745 0.275 0.835 0.74 ;
      RECT 0.745 0.275 2.59 0.365 ;
      RECT 1.565 0.865 2.255 0.955 ;
      RECT 1.07 1.045 1.97 1.135 ;
  END
END AO221X4H7R

MACRO AO222X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO222X0P5H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 1.87 0.885 1.96 1.48 ;
        RECT 1.4 1.215 1.49 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 1.79 -0.08 1.93 0.175 ;
        RECT 0.61 -0.08 0.75 0.16 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.625 0.615 1.835 0.75 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.225 0.455 1.555 0.545 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.73 0.455 1.03 0.555 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.015 0.645 1.285 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.625 0.65 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.435 0.38 0.545 ;
        RECT 0.225 0.435 0.33 0.645 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.055 0.825 2.25 0.975 ;
        RECT 2.16 0.25 2.25 0.975 ;
        RECT 2.055 0.25 2.25 0.34 ;
      LAYER MET2 ;
        RECT 2.05 0.63 2.15 1.16 ;
      LAYER VIA1 ;
        RECT 2.055 0.855 2.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.84 0.45 0.93 ;
      RECT 0.045 0.25 0.135 0.93 ;
      RECT 1.98 0.525 2.07 0.665 ;
      RECT 1.969 0.485 1.98 0.614 ;
      RECT 1.923 0.457 1.969 0.585 ;
      RECT 1.877 0.411 1.923 0.539 ;
      RECT 1.877 0.508 2.014 0.539 ;
      RECT 1.831 0.365 1.877 0.493 ;
      RECT 1.785 0.319 1.831 0.447 ;
      RECT 1.739 0.273 1.785 0.401 ;
      RECT 1.701 0.319 1.831 0.359 ;
      RECT 0.045 0.25 1.739 0.34 ;
      RECT 0.045 1.02 1.27 1.11 ;
      RECT 0.635 0.885 0.725 1.11 ;
      RECT 0.865 0.84 1.735 0.93 ;
  END
END AO222X0P5H7R

MACRO AO222X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO222X0P7H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 1.87 0.885 1.96 1.48 ;
        RECT 1.4 1.215 1.49 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 1.79 -0.08 1.93 0.175 ;
        RECT 0.61 -0.08 0.75 0.16 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.625 0.615 1.835 0.75 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.225 0.455 1.555 0.545 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.73 0.455 1.03 0.555 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.015 0.645 1.285 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.625 0.65 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.435 0.38 0.545 ;
        RECT 0.225 0.435 0.33 0.645 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.055 0.825 2.25 0.975 ;
        RECT 2.16 0.25 2.25 0.975 ;
        RECT 2.055 0.25 2.25 0.34 ;
      LAYER MET2 ;
        RECT 2.05 0.63 2.15 1.16 ;
      LAYER VIA1 ;
        RECT 2.055 0.855 2.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.84 0.45 0.93 ;
      RECT 0.045 0.25 0.135 0.93 ;
      RECT 1.98 0.525 2.07 0.665 ;
      RECT 1.969 0.485 1.98 0.614 ;
      RECT 1.923 0.457 1.969 0.585 ;
      RECT 1.877 0.411 1.923 0.539 ;
      RECT 1.877 0.508 2.014 0.539 ;
      RECT 1.831 0.365 1.877 0.493 ;
      RECT 1.785 0.319 1.831 0.447 ;
      RECT 1.739 0.273 1.785 0.401 ;
      RECT 1.701 0.319 1.831 0.359 ;
      RECT 0.045 0.25 1.739 0.34 ;
      RECT 0.045 1.02 1.27 1.11 ;
      RECT 0.635 0.885 0.725 1.11 ;
      RECT 0.865 0.84 1.735 0.93 ;
  END
END AO222X0P7H7R

MACRO AO222X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO222X1H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 1.87 0.885 1.96 1.48 ;
        RECT 1.4 1.215 1.49 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 1.79 -0.08 1.93 0.175 ;
        RECT 0.61 -0.08 0.75 0.16 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.625 0.615 1.835 0.75 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.225 0.455 1.555 0.545 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.73 0.455 1.03 0.555 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.015 0.645 1.285 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.625 0.65 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.435 0.38 0.545 ;
        RECT 0.225 0.435 0.33 0.645 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.055 0.825 2.25 0.975 ;
        RECT 2.16 0.25 2.25 0.975 ;
        RECT 2.055 0.25 2.25 0.34 ;
      LAYER MET2 ;
        RECT 2.05 0.63 2.15 1.16 ;
      LAYER VIA1 ;
        RECT 2.055 0.855 2.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.84 0.45 0.93 ;
      RECT 0.045 0.25 0.135 0.93 ;
      RECT 1.98 0.525 2.07 0.665 ;
      RECT 1.969 0.485 1.98 0.614 ;
      RECT 1.923 0.457 1.969 0.585 ;
      RECT 1.877 0.411 1.923 0.539 ;
      RECT 1.877 0.508 2.014 0.539 ;
      RECT 1.831 0.365 1.877 0.493 ;
      RECT 1.785 0.319 1.831 0.447 ;
      RECT 1.739 0.273 1.785 0.401 ;
      RECT 1.701 0.319 1.831 0.359 ;
      RECT 0.045 0.25 1.739 0.34 ;
      RECT 0.045 1.02 1.27 1.11 ;
      RECT 0.635 0.885 0.725 1.11 ;
      RECT 0.865 0.84 1.735 0.93 ;
  END
END AO222X1H7R

MACRO AO222X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO222X1P4H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 1.87 0.885 1.96 1.48 ;
        RECT 1.4 1.215 1.49 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 1.79 -0.08 1.93 0.175 ;
        RECT 0.61 -0.08 0.75 0.16 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.625 0.615 1.835 0.75 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.225 0.455 1.555 0.545 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.73 0.455 1.03 0.555 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.015 0.645 1.285 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.625 0.65 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.435 0.38 0.545 ;
        RECT 0.225 0.435 0.33 0.645 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.055 0.825 2.25 0.975 ;
        RECT 2.16 0.25 2.25 0.975 ;
        RECT 2.11 0.25 2.25 0.34 ;
      LAYER MET2 ;
        RECT 2.05 0.63 2.15 1.16 ;
      LAYER VIA1 ;
        RECT 2.055 0.855 2.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.84 0.45 0.93 ;
      RECT 0.045 0.25 0.135 0.93 ;
      RECT 1.98 0.525 2.07 0.665 ;
      RECT 1.969 0.485 1.98 0.614 ;
      RECT 1.923 0.457 1.969 0.585 ;
      RECT 1.877 0.411 1.923 0.539 ;
      RECT 1.877 0.508 2.014 0.539 ;
      RECT 1.831 0.365 1.877 0.493 ;
      RECT 1.785 0.319 1.831 0.447 ;
      RECT 1.739 0.273 1.785 0.401 ;
      RECT 1.701 0.319 1.831 0.359 ;
      RECT 0.045 0.25 1.739 0.34 ;
      RECT 0.045 1.02 1.27 1.11 ;
      RECT 0.635 0.885 0.725 1.11 ;
      RECT 0.865 0.84 1.735 0.93 ;
  END
END AO222X1P4H7R

MACRO AO222X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO222X2H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 1.835 0.88 1.925 1.48 ;
        RECT 1.365 1.215 1.455 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 1.77 -0.08 1.91 0.16 ;
        RECT 0.56 -0.08 0.7 0.16 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.595 0.64 1.82 0.76 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.305 0.455 1.605 0.545 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.715 0.455 0.98 0.555 ;
        RECT 0.715 0.455 0.855 0.585 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.645 1.235 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.625 0.605 0.745 ;
        RECT 0.47 0.51 0.605 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.43 0.375 0.545 ;
        RECT 0.225 0.43 0.335 0.635 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.055 0.825 2.215 1.145 ;
        RECT 2.125 0.355 2.215 1.145 ;
      LAYER MET2 ;
        RECT 2.05 0.63 2.15 1.16 ;
      LAYER VIA1 ;
        RECT 2.055 0.855 2.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.31 0.835 0.45 1.05 ;
      RECT 0.045 0.835 0.45 0.925 ;
      RECT 0.045 0.25 0.135 0.925 ;
      RECT 1.945 0.509 2.035 0.705 ;
      RECT 1.938 0.437 1.945 0.566 ;
      RECT 1.892 0.411 1.938 0.539 ;
      RECT 1.892 0.464 1.991 0.539 ;
      RECT 1.846 0.365 1.892 0.493 ;
      RECT 1.8 0.319 1.846 0.447 ;
      RECT 1.754 0.273 1.8 0.401 ;
      RECT 1.716 0.319 1.846 0.359 ;
      RECT 0.045 0.25 1.754 0.34 ;
      RECT 0.815 0.85 0.955 1.05 ;
      RECT 0.815 0.85 1.7 0.94 ;
      RECT 0.095 1.14 1.17 1.23 ;
      RECT 1.08 1.03 1.17 1.23 ;
      RECT 0.585 0.935 0.675 1.23 ;
      RECT 0.095 1.015 0.185 1.23 ;
      RECT 1.08 1.03 1.22 1.12 ;
      RECT 0.045 1.015 0.185 1.105 ;
  END
END AO222X2H7R

MACRO AO222X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO222X3H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 2.378 0.96 2.468 1.48 ;
        RECT 1.878 0.94 1.968 1.48 ;
        RECT 1.325 1.24 1.465 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 2.418 -0.08 2.508 0.345 ;
        RECT 1.813 -0.08 1.953 0.16 ;
        RECT 0.56 -0.08 0.7 0.16 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.625 0.61 1.825 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.39 0.455 1.48 0.6 ;
        RECT 1.225 0.455 1.48 0.545 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.74 0.455 0.975 0.545 ;
        RECT 0.74 0.455 0.83 0.625 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.645 1.235 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.42 0.625 0.645 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.43 0.375 0.545 ;
        RECT 0.225 0.43 0.33 0.64 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.103 0.835 2.258 0.925 ;
        RECT 2.168 0.255 2.258 0.925 ;
        RECT 2.025 0.255 2.258 0.345 ;
      LAYER MET2 ;
        RECT 2.05 0.18 2.15 0.56 ;
      LAYER VIA1 ;
        RECT 2.055 0.255 2.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.31 0.84 0.45 0.995 ;
      RECT 0.045 0.84 0.45 0.93 ;
      RECT 0.045 0.25 0.135 0.93 ;
      RECT 1.973 0.494 2.063 0.705 ;
      RECT 1.935 0.407 1.973 0.535 ;
      RECT 1.935 0.449 2.019 0.535 ;
      RECT 1.889 0.365 1.935 0.493 ;
      RECT 1.843 0.319 1.889 0.447 ;
      RECT 1.797 0.273 1.843 0.401 ;
      RECT 1.759 0.319 1.889 0.359 ;
      RECT 0.045 0.25 1.797 0.34 ;
      RECT 0.815 0.84 0.955 0.995 ;
      RECT 0.815 0.84 1.743 0.93 ;
      RECT 0.095 1.14 1.17 1.23 ;
      RECT 1.08 1.02 1.17 1.23 ;
      RECT 0.585 0.945 0.675 1.23 ;
      RECT 0.095 1.02 0.185 1.23 ;
      RECT 1.08 1.02 1.22 1.11 ;
      RECT 0.045 1.02 0.185 1.11 ;
  END
END AO222X3H7R

MACRO AO222X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO222X4H7R 0 0 ;
  SIZE 2.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.8 1.48 ;
        RECT 2.35 0.855 2.44 1.48 ;
        RECT 1.85 1 1.94 1.48 ;
        RECT 1.325 1.025 1.465 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.8 0.08 ;
        RECT 2.39 -0.08 2.48 0.345 ;
        RECT 1.785 -0.08 1.925 0.16 ;
        RECT 0.56 -0.08 0.7 0.16 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.623 0.595 1.803 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.39 0.455 1.48 0.65 ;
        RECT 1.225 0.455 1.48 0.545 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.74 0.455 0.975 0.545 ;
        RECT 0.74 0.455 0.83 0.675 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.645 1.235 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.625 0.65 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.455 0.375 0.545 ;
        RECT 0.225 0.455 0.315 0.695 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.115 0.395 2.255 0.485 ;
        RECT 2.055 0.825 2.215 1.145 ;
        RECT 2.115 0.395 2.215 1.145 ;
      LAYER MET2 ;
        RECT 2.05 0.63 2.15 1.16 ;
      LAYER VIA1 ;
        RECT 2.055 0.855 2.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.31 0.845 0.45 0.96 ;
      RECT 0.045 0.845 0.45 0.935 ;
      RECT 0.045 0.25 0.135 0.935 ;
      RECT 1.93 0.5 2.02 0.705 ;
      RECT 1.907 0.399 1.93 0.528 ;
      RECT 1.907 0.478 2.019 0.528 ;
      RECT 1.861 0.365 1.907 0.493 ;
      RECT 1.861 0.434 1.976 0.493 ;
      RECT 1.815 0.319 1.861 0.447 ;
      RECT 1.769 0.273 1.815 0.401 ;
      RECT 1.731 0.319 1.861 0.359 ;
      RECT 0.045 0.25 1.769 0.34 ;
      RECT 0.815 0.84 0.955 0.96 ;
      RECT 0.815 0.84 1.715 0.93 ;
      RECT 0.095 1.14 1.17 1.23 ;
      RECT 1.08 1.045 1.17 1.23 ;
      RECT 0.585 1.005 0.675 1.23 ;
      RECT 0.095 1.045 0.185 1.23 ;
      RECT 1.08 1.045 1.22 1.135 ;
      RECT 0.045 1.045 0.185 1.135 ;
  END
END AO222X4H7R

MACRO AO22X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22X0P5H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.315 0.82 1.405 1.48 ;
        RECT 0.31 1.015 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.085 -0.08 1.175 0.33 ;
        RECT 0.06 -0.08 0.2 0.315 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.425 0.235 0.575 ;
      LAYER MET2 ;
        RECT 0.05 0.23 0.15 0.76 ;
      LAYER VIA1 ;
        RECT 0.055 0.455 0.145 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.29 0.655 0.59 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.625 1.195 0.825 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.65 0.425 0.785 0.58 ;
        RECT 0.59 0.425 0.785 0.56 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.565 0.23 1.655 0.92 ;
        RECT 1.355 0.23 1.655 0.345 ;
      LAYER MET2 ;
        RECT 1.45 0.18 1.55 0.56 ;
      LAYER VIA1 ;
        RECT 1.455 0.255 1.545 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.81 0.945 0.965 1.035 ;
      RECT 0.875 0.245 0.965 1.035 ;
      RECT 1.31 0.445 1.4 0.585 ;
      RECT 0.875 0.445 1.4 0.535 ;
      RECT 0.875 0.245 0.97 0.535 ;
      RECT 0.56 0.245 0.97 0.335 ;
      RECT 0.585 1.125 1.175 1.215 ;
      RECT 1.085 0.975 1.175 1.215 ;
      RECT 0.585 0.835 0.675 1.215 ;
      RECT 0.07 0.835 0.16 1.075 ;
      RECT 0.07 0.835 0.675 0.925 ;
  END
END AO22X0P5H7R

MACRO AO22X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22X0P7H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.315 0.9 1.405 1.48 ;
        RECT 0.31 1.015 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.085 -0.08 1.175 0.33 ;
        RECT 0.06 -0.08 0.2 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.425 0.235 0.575 ;
      LAYER MET2 ;
        RECT 0.05 0.23 0.15 0.76 ;
      LAYER VIA1 ;
        RECT 0.055 0.455 0.145 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.295 0.655 0.595 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 0.62 1.185 0.82 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.67 0.425 0.775 0.58 ;
        RECT 0.58 0.425 0.775 0.55 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.565 0.255 1.655 0.968 ;
        RECT 1.355 0.255 1.655 0.345 ;
      LAYER MET2 ;
        RECT 1.45 0.18 1.55 0.56 ;
      LAYER VIA1 ;
        RECT 1.455 0.255 1.545 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.81 0.945 0.96 1.035 ;
      RECT 0.87 0.245 0.96 1.035 ;
      RECT 1.31 0.44 1.4 0.605 ;
      RECT 0.87 0.44 1.4 0.53 ;
      RECT 0.56 0.245 0.96 0.335 ;
      RECT 0.585 1.125 1.175 1.215 ;
      RECT 1.085 0.975 1.175 1.215 ;
      RECT 0.585 0.835 0.675 1.215 ;
      RECT 0.07 0.835 0.16 1.075 ;
      RECT 0.07 0.835 0.675 0.925 ;
  END
END AO22X0P7H7R

MACRO AO22X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22X1H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.3 0.9 1.39 1.48 ;
        RECT 0.295 1.015 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.07 -0.08 1.16 0.33 ;
        RECT 0.06 -0.08 0.2 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.425 0.235 0.575 ;
      LAYER MET2 ;
        RECT 0.05 0.23 0.15 0.76 ;
      LAYER VIA1 ;
        RECT 0.055 0.455 0.145 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.28 0.655 0.58 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.035 0.625 1.17 0.825 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.425 0.76 0.58 ;
        RECT 0.565 0.425 0.76 0.55 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.55 0.255 1.64 0.92 ;
        RECT 1.34 0.255 1.64 0.345 ;
      LAYER MET2 ;
        RECT 1.45 0.18 1.55 0.56 ;
      LAYER VIA1 ;
        RECT 1.455 0.255 1.545 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.795 0.945 0.945 1.035 ;
      RECT 0.855 0.245 0.945 1.035 ;
      RECT 1.295 0.445 1.385 0.605 ;
      RECT 0.855 0.445 1.385 0.535 ;
      RECT 0.545 0.245 0.945 0.335 ;
      RECT 0.57 1.125 1.16 1.215 ;
      RECT 1.07 0.975 1.16 1.215 ;
      RECT 0.57 0.835 0.66 1.215 ;
      RECT 0.07 0.835 0.16 1.075 ;
      RECT 0.07 0.835 0.66 0.925 ;
  END
END AO22X1H7R

MACRO AO22X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22X1P4H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.315 0.944 1.405 1.48 ;
        RECT 0.31 1.015 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.085 -0.08 1.175 0.33 ;
        RECT 0.06 -0.08 0.2 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.425 0.235 0.575 ;
      LAYER MET2 ;
        RECT 0.05 0.23 0.15 0.76 ;
      LAYER VIA1 ;
        RECT 0.055 0.455 0.145 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.295 0.655 0.595 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 0.625 1.185 0.825 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.685 0.425 0.775 0.607 ;
        RECT 0.58 0.425 0.775 0.545 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.565 0.255 1.655 0.92 ;
        RECT 1.355 0.255 1.655 0.345 ;
      LAYER MET2 ;
        RECT 1.45 0.18 1.55 0.56 ;
      LAYER VIA1 ;
        RECT 1.455 0.255 1.545 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.81 0.945 0.96 1.035 ;
      RECT 0.87 0.245 0.96 1.035 ;
      RECT 1.31 0.445 1.4 0.626 ;
      RECT 0.87 0.445 1.4 0.535 ;
      RECT 0.56 0.245 0.96 0.335 ;
      RECT 0.585 1.125 1.175 1.215 ;
      RECT 1.085 0.975 1.175 1.215 ;
      RECT 0.585 0.835 0.675 1.215 ;
      RECT 0.07 0.835 0.16 1.075 ;
      RECT 0.07 0.835 0.675 0.925 ;
  END
END AO22X1P4H7R

MACRO AO22X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22X2H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.315 0.855 1.405 1.48 ;
        RECT 0.31 1.015 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.615 -0.08 1.755 0.32 ;
        RECT 1.085 -0.08 1.175 0.33 ;
        RECT 0.06 -0.08 0.2 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.425 0.235 0.575 ;
      LAYER MET2 ;
        RECT 0.05 0.23 0.15 0.76 ;
      LAYER VIA1 ;
        RECT 0.055 0.455 0.145 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.295 0.655 0.595 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.75 1.192 0.885 ;
        RECT 1.055 0.62 1.145 0.885 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.577 0.425 0.78 0.56 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.56 1.025 1.745 1.175 ;
        RECT 1.56 0.523 1.655 1.175 ;
        RECT 1.542 0.499 1.652 0.55 ;
        RECT 1.496 0.453 1.606 0.518 ;
        RECT 1.45 0.421 1.56 0.472 ;
        RECT 1.423 0.389 1.542 0.436 ;
        RECT 1.377 0.343 1.496 0.399 ;
        RECT 1.331 0.22 1.45 0.353 ;
        RECT 1.3 0.22 1.45 0.33 ;
      LAYER MET2 ;
        RECT 1.65 0.84 1.75 1.22 ;
      LAYER VIA1 ;
        RECT 1.655 1.055 1.745 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.81 0.945 0.96 1.035 ;
      RECT 0.87 0.215 0.96 1.035 ;
      RECT 1.265 0.463 1.355 0.626 ;
      RECT 0.87 0.44 1.309 0.53 ;
      RECT 0.56 0.215 0.96 0.305 ;
      RECT 0.585 1.125 1.175 1.215 ;
      RECT 1.085 0.975 1.175 1.215 ;
      RECT 0.585 0.835 0.675 1.215 ;
      RECT 0.07 0.835 0.16 1.075 ;
      RECT 0.07 0.835 0.675 0.925 ;
  END
END AO22X2H7R

MACRO AO22X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22X3H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.815 0.915 1.905 1.48 ;
        RECT 1.315 0.915 1.405 1.48 ;
        RECT 0.31 1.015 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.63 -0.08 1.72 0.345 ;
        RECT 1.085 -0.08 1.175 0.33 ;
        RECT 0.06 -0.08 0.2 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.425 0.26 0.555 ;
        RECT 0.055 0.425 0.145 0.575 ;
      LAYER MET2 ;
        RECT 0.05 0.23 0.15 0.76 ;
      LAYER VIA1 ;
        RECT 0.055 0.455 0.145 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.29 0.655 0.59 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 0.625 1.18 0.857 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.64 0.425 0.78 0.58 ;
        RECT 0.595 0.425 0.78 0.545 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.655 0.591 1.745 0.825 ;
        RECT 1.655 0.559 1.726 0.857 ;
        RECT 1.54 0.79 1.68 0.88 ;
        RECT 1.655 0.523 1.68 0.88 ;
        RECT 1.642 0.783 1.745 0.825 ;
        RECT 1.654 0.51 1.655 0.639 ;
        RECT 1.608 0.487 1.654 0.615 ;
        RECT 1.516 0.441 1.608 0.523 ;
        RECT 1.562 0.441 1.608 0.569 ;
        RECT 1.47 0.395 1.562 0.477 ;
        RECT 1.426 0.349 1.516 0.432 ;
        RECT 1.38 0.22 1.47 0.387 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.81 0.885 0.96 0.975 ;
      RECT 0.87 0.245 0.96 0.975 ;
      RECT 1.28 0.503 1.37 0.686 ;
      RECT 1.261 0.503 1.37 0.545 ;
      RECT 0.87 0.445 1.299 0.535 ;
      RECT 0.87 0.468 1.345 0.535 ;
      RECT 0.56 0.245 0.96 0.335 ;
      RECT 0.585 1.065 1.175 1.155 ;
      RECT 1.085 0.975 1.175 1.155 ;
      RECT 0.585 0.835 0.675 1.155 ;
      RECT 0.07 0.835 0.16 1.015 ;
      RECT 0.07 0.835 0.675 0.925 ;
  END
END AO22X3H7R

MACRO AO22X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22X4H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.805 1.035 1.945 1.48 ;
        RECT 1.33 0.81 1.42 1.48 ;
        RECT 0.31 1.095 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.62 -0.08 1.76 0.235 ;
        RECT 1.085 -0.08 1.175 0.365 ;
        RECT 0.085 -0.08 0.175 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.38 0.625 0.56 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.685 1.145 0.995 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.425 0.775 0.66 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.555 0.855 2 0.945 ;
        RECT 1.91 0.275 2 0.945 ;
        RECT 1.38 0.325 2 0.415 ;
        RECT 1.38 0.25 1.47 0.415 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.81 0.905 0.96 0.995 ;
      RECT 0.87 0.245 0.96 0.995 ;
      RECT 0.87 0.505 1.625 0.595 ;
      RECT 0.56 0.245 0.96 0.335 ;
      RECT 0.585 1.085 1.2 1.175 ;
      RECT 0.585 0.915 0.675 1.175 ;
      RECT 0.07 0.915 0.16 1.055 ;
      RECT 0.07 0.915 0.675 1.005 ;
  END
END AO22X4H7R

MACRO AO22X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22X6H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 1.805 1.035 1.945 1.48 ;
        RECT 1.33 0.81 1.42 1.48 ;
        RECT 0.31 1.095 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 2.18 -0.08 2.27 0.37 ;
        RECT 1.635 -0.08 1.775 0.235 ;
        RECT 1.085 -0.08 1.175 0.365 ;
        RECT 0.085 -0.08 0.175 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.605 0.56 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.685 1.155 0.975 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.425 0.775 0.685 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.08 0.79 2.17 1.13 ;
        RECT 2 0.325 2.09 0.945 ;
        RECT 1.58 0.855 2.17 0.945 ;
        RECT 1.37 0.325 2.09 0.415 ;
        RECT 1.58 0.79 1.67 1.13 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.81 0.905 0.96 0.995 ;
      RECT 0.87 0.245 0.96 0.995 ;
      RECT 1.315 0.555 1.855 0.645 ;
      RECT 0.87 0.505 1.4 0.595 ;
      RECT 0.56 0.245 0.96 0.335 ;
      RECT 0.585 1.085 1.2 1.175 ;
      RECT 0.585 0.915 0.675 1.175 ;
      RECT 0.07 0.915 0.16 1.055 ;
      RECT 0.07 0.915 0.675 1.005 ;
  END
END AO22X6H7R

MACRO AO31X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO31X0P5H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.39 1.015 1.48 1.48 ;
        RECT 0.56 1.225 0.7 1.48 ;
        RECT 0.07 1.015 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.075 -0.08 1.215 0.16 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.26 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.405 0.785 0.575 0.945 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.54 0.455 0.81 0.555 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.655 1.095 0.755 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.64 0.225 1.745 1.175 ;
      LAYER MET2 ;
        RECT 1.65 0.84 1.75 1.22 ;
      LAYER VIA1 ;
        RECT 1.655 1.055 1.745 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.075 1.04 1.3 1.13 ;
      RECT 1.21 0.25 1.3 1.13 ;
      RECT 1.21 0.58 1.55 0.67 ;
      RECT 0.795 0.25 1.3 0.34 ;
      RECT 0.295 1.045 0.965 1.135 ;
  END
END AO31X0P5H7R

MACRO AO31X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO31X0P7H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.39 1.035 1.48 1.48 ;
        RECT 0.56 1.215 0.7 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.39 -0.08 1.48 0.365 ;
        RECT 1.08 -0.08 1.17 0.365 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.405 0.785 0.575 0.945 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.54 0.455 0.81 0.555 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.655 1.05 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.64 0.225 1.745 1.103 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.56 ;
      LAYER VIA1 ;
        RECT 1.655 0.255 1.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.075 1.02 1.23 1.11 ;
      RECT 1.14 0.475 1.23 1.11 ;
      RECT 1.14 0.58 1.55 0.67 ;
      RECT 0.9 0.475 1.23 0.565 ;
      RECT 0.9 0.26 0.99 0.565 ;
      RECT 0.795 0.26 0.99 0.35 ;
      RECT 0.295 1.035 0.965 1.125 ;
  END
END AO31X0P7H7R

MACRO AO31X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO31X1H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.39 1.015 1.48 1.48 ;
        RECT 0.56 1.225 0.7 1.48 ;
        RECT 0.07 1.015 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.39 -0.08 1.48 0.35 ;
        RECT 1.09 -0.08 1.18 0.35 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.26 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.395 0.795 0.575 0.945 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 0.455 0.82 0.555 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.655 1.095 0.755 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.64 0.225 1.745 1.175 ;
      LAYER MET2 ;
        RECT 1.65 0.84 1.75 1.22 ;
      LAYER VIA1 ;
        RECT 1.655 1.055 1.745 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.075 1.04 1.3 1.13 ;
      RECT 1.21 0.475 1.3 1.13 ;
      RECT 1.21 0.58 1.55 0.67 ;
      RECT 0.91 0.475 1.3 0.565 ;
      RECT 0.91 0.25 1 0.565 ;
      RECT 0.795 0.25 1 0.34 ;
      RECT 0.295 1.045 0.965 1.135 ;
  END
END AO31X1H7R

MACRO AO31X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO31X1P4H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.39 1.035 1.48 1.48 ;
        RECT 0.56 1.215 0.7 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.39 -0.08 1.48 0.365 ;
        RECT 1.09 -0.08 1.18 0.365 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.26 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.395 0.795 0.575 0.945 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 0.455 0.82 0.555 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.655 1.05 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.64 0.225 1.745 1.011 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.56 ;
      LAYER VIA1 ;
        RECT 1.655 0.255 1.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.075 1.02 1.23 1.11 ;
      RECT 1.14 0.475 1.23 1.11 ;
      RECT 1.14 0.58 1.55 0.67 ;
      RECT 0.91 0.475 1.23 0.565 ;
      RECT 0.91 0.25 1 0.565 ;
      RECT 0.795 0.25 1 0.34 ;
      RECT 0.295 1.035 0.965 1.125 ;
  END
END AO31X1P4H7R

MACRO AO31X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO31X2H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.61 1.02 1.7 1.48 ;
        RECT 1.11 1.045 1.2 1.48 ;
        RECT 0.57 1.225 0.71 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.595 -0.08 1.685 0.38 ;
        RECT 1.085 -0.08 1.175 0.365 ;
        RECT 0.045 -0.08 0.185 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.985 0.605 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.735 0.255 0.825 0.59 ;
        RECT 0.625 0.255 0.825 0.345 ;
      LAYER MET2 ;
        RECT 0.65 0.18 0.75 0.56 ;
      LAYER VIA1 ;
        RECT 0.655 0.255 0.745 0.345 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.48 0.455 0.575 0.69 ;
        RECT 0.425 0.455 0.575 0.545 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.655 0.375 0.75 ;
        RECT 0.225 0.52 0.32 0.75 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.415 0.655 1.575 0.745 ;
        RECT 1.335 1.045 1.505 1.135 ;
        RECT 1.415 0.265 1.505 1.135 ;
        RECT 1.31 0.265 1.505 0.355 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.865 0.16 1.16 ;
      RECT 0.045 0.865 1.325 0.955 ;
      RECT 1.235 0.575 1.325 0.955 ;
      RECT 0.045 0.265 0.135 1.16 ;
      RECT 0.045 0.265 0.45 0.355 ;
      RECT 0.295 1.045 0.975 1.135 ;
  END
END AO31X2H7R

MACRO AO31X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO31X3H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.61 1.03 1.7 1.48 ;
        RECT 1.11 1.045 1.2 1.48 ;
        RECT 0.57 1.225 0.71 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.595 -0.08 1.685 0.375 ;
        RECT 1.085 -0.08 1.175 0.36 ;
        RECT 0.045 -0.08 0.185 0.225 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.625 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.625 0.835 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.425 0.555 0.695 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.575 0.36 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.415 0.625 1.545 0.775 ;
        RECT 1.335 1.045 1.505 1.135 ;
        RECT 1.415 0.35 1.505 1.135 ;
        RECT 1.31 0.35 1.505 0.44 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.865 0.16 1.07 ;
      RECT 0.045 0.865 1.325 0.955 ;
      RECT 1.235 0.685 1.325 0.955 ;
      RECT 0.045 0.473 0.135 1.07 ;
      RECT 0.091 0.428 0.181 0.511 ;
      RECT 0.135 0.383 0.227 0.465 ;
      RECT 0.135 0.383 0.273 0.419 ;
      RECT 0.181 0.337 0.296 0.385 ;
      RECT 0.227 0.291 0.334 0.354 ;
      RECT 0.273 0.256 0.296 0.385 ;
      RECT 0.296 0.245 0.45 0.335 ;
      RECT 0.295 1.045 0.975 1.135 ;
  END
END AO31X3H7R

MACRO AO31X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO31X4H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.66 1.055 1.75 1.48 ;
        RECT 1.16 1.045 1.25 1.48 ;
        RECT 0.62 1.225 0.76 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.615 -0.08 1.705 0.345 ;
        RECT 1.115 -0.08 1.205 0.33 ;
        RECT 0.07 -0.08 0.16 0.245 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.015 0.595 1.165 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.625 0.835 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.425 0.565 0.675 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.245 0.55 0.365 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.385 1.045 1.545 1.135 ;
        RECT 1.455 0.526 1.545 1.135 ;
        RECT 1.411 0.481 1.501 0.564 ;
        RECT 1.365 0.355 1.455 0.519 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.065 0.865 0.21 1.01 ;
      RECT 0.065 0.865 1.355 0.955 ;
      RECT 1.265 0.615 1.355 0.955 ;
      RECT 0.065 0.448 0.155 1.01 ;
      RECT 0.111 0.403 0.201 0.486 ;
      RECT 0.155 0.358 0.247 0.44 ;
      RECT 0.201 0.312 0.291 0.395 ;
      RECT 0.201 0.312 0.329 0.354 ;
      RECT 0.291 0.245 0.5 0.335 ;
      RECT 0.247 0.267 0.5 0.335 ;
      RECT 0.345 1.045 1.025 1.135 ;
  END
END AO31X4H7R

MACRO AOA211X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOA211X0P5H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.29 1.05 1.38 1.48 ;
        RECT 0.31 1.075 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.34 -0.08 1.43 0.365 ;
        RECT 0.535 -0.08 0.675 0.16 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.26 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.405 0.655 0.585 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.525 0.435 0.795 0.545 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.84 0.625 1.02 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.59 0.225 1.745 0.375 ;
        RECT 1.515 1.02 1.68 1.11 ;
        RECT 1.59 0.225 1.68 1.11 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.56 ;
      LAYER VIA1 ;
        RECT 1.655 0.255 1.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.825 1.005 1.2 1.095 ;
      RECT 1.11 0.225 1.2 1.095 ;
      RECT 1.11 0.58 1.5 0.67 ;
      RECT 0.575 1.04 0.715 1.13 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 0.095 0.895 0.185 1.13 ;
      RECT 0.575 0.895 0.665 1.13 ;
      RECT 0.095 0.895 0.665 0.985 ;
      RECT 0.045 0.25 0.975 0.34 ;
  END
END AOA211X0P5H7R

MACRO AOA211X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOA211X0P7H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.29 1.05 1.38 1.48 ;
        RECT 0.31 1.075 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.34 -0.08 1.43 0.365 ;
        RECT 0.545 -0.08 0.685 0.16 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.26 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.405 0.655 0.585 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.525 0.435 0.795 0.545 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.84 0.625 1.02 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.59 0.225 1.745 0.375 ;
        RECT 1.515 0.99 1.68 1.08 ;
        RECT 1.59 0.225 1.68 1.08 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.56 ;
      LAYER VIA1 ;
        RECT 1.655 0.255 1.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.825 1.005 1.2 1.095 ;
      RECT 1.11 0.225 1.2 1.095 ;
      RECT 1.11 0.58 1.5 0.67 ;
      RECT 0.575 1.04 0.715 1.13 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 0.095 0.895 0.185 1.13 ;
      RECT 0.575 0.895 0.665 1.13 ;
      RECT 0.095 0.895 0.665 0.985 ;
      RECT 0.045 0.25 0.975 0.34 ;
  END
END AOA211X0P7H7R

MACRO AOA211X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOA211X1H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.29 1.05 1.38 1.48 ;
        RECT 0.31 1.075 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.34 -0.08 1.43 0.365 ;
        RECT 0.545 -0.08 0.685 0.16 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.26 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.405 0.655 0.585 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.525 0.435 0.795 0.545 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.84 0.625 1.02 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.59 0.225 1.745 0.375 ;
        RECT 1.515 0.94 1.68 1.03 ;
        RECT 1.59 0.225 1.68 1.03 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.56 ;
      LAYER VIA1 ;
        RECT 1.655 0.255 1.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.825 1.005 1.2 1.095 ;
      RECT 1.11 0.225 1.2 1.095 ;
      RECT 1.11 0.58 1.5 0.67 ;
      RECT 0.575 1.04 0.715 1.13 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 0.095 0.895 0.185 1.13 ;
      RECT 0.575 0.895 0.665 1.13 ;
      RECT 0.095 0.895 0.665 0.985 ;
      RECT 0.045 0.25 0.975 0.34 ;
  END
END AOA211X1H7R

MACRO AOA211X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOA211X1P4H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.29 1.05 1.38 1.48 ;
        RECT 0.31 1.075 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.34 -0.08 1.43 0.355 ;
        RECT 0.545 -0.08 0.685 0.16 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.26 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.405 0.655 0.585 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.525 0.435 0.795 0.545 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.84 0.625 1.02 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.825 1.68 0.975 ;
        RECT 1.59 0.31 1.68 0.975 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.825 1.005 1.2 1.095 ;
      RECT 1.11 0.225 1.2 1.095 ;
      RECT 1.11 0.58 1.5 0.67 ;
      RECT 0.575 1.04 0.715 1.13 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 0.095 0.895 0.185 1.13 ;
      RECT 0.575 0.895 0.665 1.13 ;
      RECT 0.095 0.895 0.665 0.985 ;
      RECT 0.045 0.25 0.975 0.34 ;
  END
END AOA211X1P4H7R

MACRO AOA211X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOA211X2H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.29 1.05 1.38 1.48 ;
        RECT 0.31 1.225 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.34 -0.08 1.43 0.345 ;
        RECT 0.555 -0.08 0.695 0.16 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.26 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.405 0.795 0.585 0.945 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.525 0.445 0.795 0.545 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.84 0.625 1.02 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.59 0.825 1.745 0.975 ;
        RECT 1.59 0.34 1.68 0.975 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.825 1.005 1.2 1.095 ;
      RECT 1.11 0.225 1.2 1.095 ;
      RECT 1.11 0.59 1.5 0.68 ;
      RECT 0.045 0.25 0.975 0.34 ;
      RECT 0.045 1.04 0.715 1.13 ;
  END
END AOA211X2H7R

MACRO AOA211X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOA211X3H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.835 1.035 1.925 1.48 ;
        RECT 1.33 1.05 1.42 1.48 ;
        RECT 0.31 1.225 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.83 -0.08 1.92 0.355 ;
        RECT 1.33 -0.08 1.42 0.355 ;
        RECT 0.52 -0.08 0.66 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.26 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.765 0.575 0.945 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.45 0.805 0.6 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.855 1.05 0.945 ;
        RECT 0.96 0.75 1.05 0.945 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.58 0.825 1.745 1.025 ;
        RECT 1.58 0.305 1.67 1.025 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.825 1.04 1.23 1.13 ;
      RECT 1.14 0.58 1.23 1.13 ;
      RECT 1.14 0.58 1.49 0.67 ;
      RECT 1.106 0.565 1.226 0.605 ;
      RECT 1.06 0.275 1.15 0.565 ;
      RECT 1.06 0.527 1.196 0.565 ;
      RECT 0.045 0.265 0.925 0.355 ;
      RECT 0.045 1.04 0.715 1.13 ;
  END
END AOA211X3H7R

MACRO AOA211X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOA211X4H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 1.85 1.055 1.94 1.48 ;
        RECT 1.35 1.05 1.44 1.48 ;
        RECT 0.31 1.075 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 1.89 -0.08 1.98 0.345 ;
        RECT 1.39 -0.08 1.48 0.345 ;
        RECT 0.57 -0.08 0.71 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.26 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.395 0.655 0.575 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.75 0.455 0.84 0.66 ;
        RECT 0.625 0.455 0.84 0.545 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.855 1.08 0.945 ;
        RECT 0.99 0.665 1.08 0.945 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.575 0.835 1.745 0.925 ;
        RECT 1.64 0.37 1.745 0.925 ;
      LAYER MET2 ;
        RECT 1.65 0.23 1.75 0.76 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.825 1.04 1.26 1.13 ;
      RECT 1.17 0.31 1.26 1.13 ;
      RECT 1.17 0.58 1.49 0.67 ;
      RECT 1.14 0.31 1.26 0.45 ;
      RECT 0.045 0.895 0.185 1.015 ;
      RECT 0.045 0.895 0.715 0.985 ;
      RECT 0.045 0.265 1.025 0.355 ;
  END
END AOA211X4H7R

MACRO AOAI211X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOAI211X0P5H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.16 1.035 1.25 1.48 ;
        RECT 0.31 1.075 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.545 -0.08 0.685 0.16 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.26 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.405 0.655 0.585 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.525 0.435 0.795 0.545 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.84 0.625 1.02 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.11 0.225 1.345 0.375 ;
        RECT 1.11 0.225 1.2 0.886 ;
        RECT 1.015 0.898 1.11 0.956 ;
        RECT 1.061 0.852 1.156 0.931 ;
        RECT 1.107 0.827 1.11 0.956 ;
        RECT 0.969 0.944 1.107 0.98 ;
        RECT 0.931 0.986 1.061 1.026 ;
        RECT 0.969 0.944 1.061 1.026 ;
        RECT 0.825 1.005 1.015 1.072 ;
        RECT 0.825 1.005 0.969 1.095 ;
      LAYER MET2 ;
        RECT 1.25 0.18 1.35 0.56 ;
      LAYER VIA1 ;
        RECT 1.255 0.255 1.345 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.575 1.04 0.715 1.13 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 0.095 0.895 0.185 1.13 ;
      RECT 0.575 0.895 0.665 1.13 ;
      RECT 0.095 0.895 0.665 0.985 ;
      RECT 0.045 0.25 0.975 0.34 ;
  END
END AOAI211X0P5H7R

MACRO AOAI211X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOAI211X0P7H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.155 1.035 1.245 1.48 ;
        RECT 0.31 1.075 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.545 -0.08 0.685 0.16 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.26 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.395 0.655 0.62 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.525 0.445 0.795 0.55 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.78 0.645 1.05 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.275 1.345 0.736 ;
        RECT 1.18 0.728 1.301 0.781 ;
        RECT 1.226 0.69 1.255 0.819 ;
        RECT 1.085 0.275 1.345 0.365 ;
        RECT 1.134 0.774 1.226 0.856 ;
        RECT 1.088 0.82 1.18 0.902 ;
        RECT 1.042 0.866 1.134 0.948 ;
        RECT 0.958 0.954 1.088 0.994 ;
        RECT 0.996 0.912 1.088 0.994 ;
        RECT 0.825 0.973 1.042 1.04 ;
        RECT 0.825 0.973 0.996 1.063 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.575 0.988 0.715 1.078 ;
      RECT 0.045 0.988 0.185 1.078 ;
      RECT 0.095 0.865 0.185 1.078 ;
      RECT 0.575 0.865 0.665 1.078 ;
      RECT 0.095 0.865 0.665 0.955 ;
      RECT 0.045 0.25 0.975 0.34 ;
  END
END AOAI211X0P7H7R

MACRO AOAI211X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOAI211X1H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.165 1.035 1.255 1.48 ;
        RECT 0.31 1.105 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.535 -0.08 0.675 0.16 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.26 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.655 0.575 0.835 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.61 0.455 0.81 0.545 ;
        RECT 0.675 0.455 0.765 0.645 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.625 1.035 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.31 1.345 0.746 ;
        RECT 1.146 0.772 1.255 0.823 ;
        RECT 1.192 0.726 1.301 0.791 ;
        RECT 1.238 0.694 1.255 0.823 ;
        RECT 1.085 0.31 1.345 0.4 ;
        RECT 1.1 0.818 1.238 0.854 ;
        RECT 1.1 0.818 1.192 0.9 ;
        RECT 1.016 0.906 1.146 0.946 ;
        RECT 1.054 0.864 1.146 0.946 ;
        RECT 0.825 0.925 1.1 0.992 ;
        RECT 0.825 0.925 1.054 1.015 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.925 0.185 1.045 ;
      RECT 0.045 0.925 0.715 1.015 ;
      RECT 0.045 0.25 0.975 0.34 ;
  END
END AOAI211X1H7R

MACRO AOAI211X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOAI211X1P4H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.115 1.075 1.255 1.48 ;
        RECT 0.295 1.075 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.585 -0.08 0.725 0.16 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.26 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.375 0.655 0.575 0.79 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.755 0.455 0.845 0.625 ;
        RECT 0.625 0.455 0.845 0.545 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.995 0.595 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.325 1.345 0.857 ;
        RECT 1.167 0.866 1.301 0.902 ;
        RECT 1.251 0.799 1.255 0.927 ;
        RECT 1.165 0.325 1.345 0.415 ;
        RECT 0.865 0.885 1.251 0.952 ;
        RECT 1.205 0.824 1.301 0.902 ;
        RECT 0.865 0.885 1.205 0.975 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.895 0.185 1.015 ;
      RECT 0.045 0.895 0.695 0.985 ;
      RECT 0.045 0.25 1.055 0.34 ;
  END
END AOAI211X1P4H7R

MACRO AOAI211X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOAI211X2H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.332 1.055 1.422 1.48 ;
        RECT 0.532 1.07 0.622 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 0.797 -0.08 0.937 0.185 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.645 0.495 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.585 0.64 0.785 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.962 0.455 1.052 0.69 ;
        RECT 0.825 0.455 1.052 0.545 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.195 0.595 1.345 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.057 0.865 1.545 0.955 ;
        RECT 1.455 0.34 1.545 0.955 ;
        RECT 1.377 0.34 1.545 0.43 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.257 0.275 1.267 0.365 ;
      RECT 0.257 0.89 0.897 0.98 ;
  END
END AOAI211X2H7R

MACRO AOAI211X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOAI211X3H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 2.025 1.095 2.165 1.48 ;
        RECT 1.045 1.08 1.185 1.48 ;
        RECT 0.545 1.08 0.685 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 1.555 -0.08 1.695 0.335 ;
        RECT 0.295 -0.08 0.435 0.335 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.695 0.655 1.035 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.165 0.655 0.505 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.425 0.655 1.765 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.925 0.655 2.265 0.745 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.8 0.915 2.545 1.005 ;
        RECT 2.455 0.465 2.545 1.005 ;
        RECT 2.07 0.465 2.545 0.555 ;
        RECT 2.3 0.915 2.39 1.06 ;
        RECT 2.07 0.35 2.21 0.555 ;
        RECT 1.275 1.11 1.89 1.2 ;
        RECT 1.8 0.915 1.89 1.2 ;
        RECT 1.275 1.08 1.415 1.2 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.81 0.44 1.92 0.53 ;
      RECT 1.83 0.17 1.92 0.53 ;
      RECT 1.33 0.28 1.42 0.53 ;
      RECT 0.81 0.35 0.95 0.53 ;
      RECT 2.36 0.17 2.45 0.375 ;
      RECT 1.83 0.17 2.45 0.26 ;
      RECT 0.82 0.9 0.91 1.045 ;
      RECT 0.32 0.9 0.41 1.045 ;
      RECT 1.525 0.9 1.665 1.02 ;
      RECT 0.32 0.9 1.665 0.99 ;
      RECT 0.07 0.425 0.66 0.515 ;
      RECT 0.57 0.17 0.66 0.515 ;
      RECT 0.07 0.28 0.16 0.515 ;
      RECT 1.075 0.17 1.215 0.35 ;
      RECT 0.57 0.17 1.215 0.26 ;
  END
END AOAI211X3H7R

MACRO AOAI211X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOAI211X4H7R 0 0 ;
  SIZE 3 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3 1.48 ;
        RECT 2.262 1.07 2.352 1.48 ;
        RECT 1.257 1.08 1.397 1.48 ;
        RECT 0.782 1.07 0.872 1.48 ;
        RECT 0.282 1.055 0.372 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3 0.08 ;
        RECT 1.767 -0.08 1.907 0.305 ;
        RECT 0.507 -0.08 0.647 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.907 0.655 1.247 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.377 0.655 0.717 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.637 0.655 1.977 0.745 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.137 0.655 2.477 0.745 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.012 0.855 2.657 0.945 ;
        RECT 2.567 0.553 2.657 0.945 ;
        RECT 2.523 0.508 2.613 0.591 ;
        RECT 2.477 0.463 2.567 0.546 ;
        RECT 2.282 0.418 2.523 0.485 ;
        RECT 2.282 0.395 2.477 0.485 ;
        RECT 2.439 0.463 2.567 0.504 ;
        RECT 1.487 1.065 2.102 1.155 ;
        RECT 2.012 0.855 2.102 1.155 ;
      LAYER MET2 ;
        RECT 2.45 0.625 2.55 1.16 ;
      LAYER VIA1 ;
        RECT 2.455 0.855 2.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.022 0.41 2.132 0.507 ;
      RECT 2.042 0.215 2.132 0.507 ;
      RECT 1.517 0.38 1.657 0.507 ;
      RECT 1.022 0.395 1.162 0.507 ;
      RECT 2.572 0.215 2.662 0.355 ;
      RECT 2.042 0.215 2.662 0.305 ;
      RECT 0.282 0.395 0.872 0.485 ;
      RECT 0.782 0.215 0.872 0.485 ;
      RECT 0.282 0.28 0.372 0.485 ;
      RECT 1.287 0.215 1.427 0.32 ;
      RECT 0.782 0.215 1.427 0.305 ;
      RECT 0.507 0.885 1.877 0.975 ;
  END
END AOAI211X4H7R

MACRO AOI211X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211X0P5H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.015 -0.08 1.155 0.32 ;
        RECT 0.505 -0.08 0.645 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.6 0.545 0.8 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.905 0.645 1.175 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.25 1.15 0.785 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.68 0.855 0.975 0.945 ;
        RECT 0.68 0.805 0.77 0.945 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.015 1.055 1.355 1.145 ;
        RECT 1.265 0.41 1.355 1.145 ;
        RECT 0.07 0.41 1.355 0.5 ;
        RECT 0.78 0.22 0.87 0.5 ;
        RECT 0.07 0.205 0.16 0.5 ;
      LAYER MET2 ;
        RECT 1.05 1.015 1.15 1.22 ;
      LAYER VIA1 ;
        RECT 1.055 1.055 1.145 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.57 1.034 0.66 1.2 ;
      RECT 0.07 0.915 0.16 1.155 ;
      RECT 0.565 0.963 0.57 1.092 ;
      RECT 0.519 0.938 0.565 1.066 ;
      RECT 0.519 0.989 0.616 1.066 ;
      RECT 0.481 0.989 0.616 1.024 ;
      RECT 0.07 0.915 0.519 1.005 ;
  END
END AOI211X0P5H7R

MACRO AOI211X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211X0P7H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.025 -0.08 1.165 0.32 ;
        RECT 0.505 -0.08 0.645 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.6 0.545 0.8 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.905 0.645 1.175 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.25 1.15 0.785 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.736 0.855 0.975 0.945 ;
        RECT 0.69 0.755 0.78 0.922 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 1.055 1.355 1.145 ;
        RECT 1.265 0.41 1.355 1.145 ;
        RECT 0.07 0.41 1.355 0.5 ;
        RECT 0.78 0.245 0.87 0.5 ;
        RECT 0.07 0.23 0.16 0.5 ;
      LAYER MET2 ;
        RECT 1.05 1.015 1.15 1.22 ;
      LAYER VIA1 ;
        RECT 1.055 1.055 1.145 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.57 0.981 0.66 1.145 ;
      RECT 0.07 0.915 0.16 1.123 ;
      RECT 0.536 0.981 0.66 1.022 ;
      RECT 0.07 0.915 0.574 1.005 ;
      RECT 0.07 0.938 0.62 1.005 ;
  END
END AOI211X0P7H7R

MACRO AOI211X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211X1H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.035 -0.08 1.175 0.32 ;
        RECT 0.505 -0.08 0.645 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.6 0.545 0.8 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.045 0.625 1.145 0.785 ;
        RECT 0.905 0.625 1.145 0.765 ;
      LAYER MET2 ;
        RECT 1.05 0.25 1.15 0.785 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.716 0.855 0.98 0.945 ;
        RECT 0.68 0.725 0.77 0.927 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 1.055 1.325 1.145 ;
        RECT 1.235 0.41 1.325 1.145 ;
        RECT 0.07 0.41 1.325 0.5 ;
        RECT 0.78 0.28 0.87 0.5 ;
        RECT 0.07 0.265 0.16 0.5 ;
      LAYER MET2 ;
        RECT 1.05 1.015 1.15 1.22 ;
      LAYER VIA1 ;
        RECT 1.055 1.055 1.145 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.57 1.034 0.66 1.2 ;
      RECT 0.07 0.915 0.16 1.17 ;
      RECT 0.565 0.963 0.57 1.092 ;
      RECT 0.519 0.938 0.565 1.066 ;
      RECT 0.519 0.989 0.616 1.066 ;
      RECT 0.481 0.989 0.616 1.024 ;
      RECT 0.07 0.915 0.519 1.005 ;
  END
END AOI211X1H7R

MACRO AOI211X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211X1P4H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.02 -0.08 1.16 0.32 ;
        RECT 0.505 -0.08 0.645 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.6 0.545 0.8 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.905 0.645 1.175 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.25 1.15 0.785 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.801 0.855 0.98 0.945 ;
        RECT 0.726 0.836 0.839 0.892 ;
        RECT 0.68 0.801 0.801 0.847 ;
        RECT 0.77 0.855 0.98 0.93 ;
        RECT 0.68 0.681 0.77 0.847 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.005 1.055 1.355 1.145 ;
        RECT 1.265 0.41 1.355 1.145 ;
        RECT 0.07 0.41 1.355 0.5 ;
        RECT 0.78 0.315 0.87 0.5 ;
        RECT 0.07 0.3 0.16 0.5 ;
      LAYER MET2 ;
        RECT 1.05 1.015 1.15 1.22 ;
      LAYER VIA1 ;
        RECT 1.055 1.055 1.145 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.585 0.933 0.675 1.091 ;
      RECT 0.07 0.915 0.16 1.055 ;
      RECT 0.07 0.915 0.639 1.005 ;
  END
END AOI211X1P4H7R

MACRO AOI211X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211X2H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 0.573 1.07 0.663 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.258 -0.08 1.398 0.305 ;
        RECT 0.758 -0.08 0.898 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.623 0.625 0.803 0.775 ;
      LAYER MET2 ;
        RECT 0.689 0.43 0.789 0.96 ;
      LAYER VIA1 ;
        RECT 0.694 0.655 0.784 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.249 0.625 0.474 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.294 0.625 1.384 0.775 ;
        RECT 1.144 0.625 1.384 0.715 ;
      LAYER MET2 ;
        RECT 1.289 0.255 1.389 0.785 ;
      LAYER VIA1 ;
        RECT 1.294 0.655 1.384 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.064 0.855 1.214 0.945 ;
        RECT 0.979 0.836 1.102 0.882 ;
        RECT 0.933 0.796 1.064 0.837 ;
        RECT 1.023 0.855 1.214 0.925 ;
        RECT 0.933 0.615 1.023 0.837 ;
      LAYER MET2 ;
        RECT 1.089 0.63 1.189 1.16 ;
      LAYER VIA1 ;
        RECT 1.094 0.855 1.184 0.945 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.258 1.055 1.564 1.145 ;
        RECT 1.474 0.395 1.564 1.145 ;
        RECT 0.323 0.395 1.564 0.485 ;
        RECT 0.323 0.295 0.413 0.485 ;
      LAYER MET2 ;
        RECT 1.289 1.015 1.389 1.22 ;
      LAYER VIA1 ;
        RECT 1.294 1.055 1.384 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.823 0.903 0.913 1.07 ;
      RECT 0.298 0.88 0.867 0.97 ;
  END
END AOI211X2H7R

MACRO AOI211X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211X3H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 0.84 1.225 0.98 1.48 ;
        RECT 0.31 1.225 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 2.15 -0.08 2.24 0.365 ;
        RECT 1.61 -0.08 1.75 0.185 ;
        RECT 1.005 -0.08 1.145 0.305 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.22 0.855 1.02 0.945 ;
        RECT 0.93 0.69 1.02 0.945 ;
        RECT 0.22 0.69 0.31 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.655 0.785 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.695 0.455 1.835 0.6 ;
        RECT 1.62 0.455 1.835 0.545 ;
      LAYER MET2 ;
        RECT 1.65 0.23 1.75 0.76 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.577 0.695 2.095 0.785 ;
        RECT 1.29 0.676 1.615 0.745 ;
        RECT 1.29 0.657 1.577 0.745 ;
        RECT 1.575 0.695 2.095 0.783 ;
        RECT 1.29 0.655 1.575 0.745 ;
        RECT 1.537 0.695 2.095 0.764 ;
        RECT 1.29 0.605 1.38 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.33 0.275 2.015 0.365 ;
        RECT 1.456 0.91 1.735 1 ;
        RECT 1.11 0.891 1.494 0.945 ;
        RECT 1.11 0.863 1.456 0.945 ;
        RECT 1.439 0.91 1.735 0.992 ;
        RECT 1.11 0.855 1.439 0.945 ;
        RECT 1.401 0.91 1.735 0.964 ;
        RECT 0.55 0.395 1.42 0.485 ;
        RECT 1.33 0.275 1.42 0.485 ;
        RECT 1.11 0.395 1.2 0.945 ;
        RECT 0.55 0.295 0.64 0.485 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.352 1.09 1.84 1.18 ;
      RECT 1.345 1.048 1.352 1.177 ;
      RECT 1.345 1.09 1.87 1.165 ;
      RECT 1.307 1.09 1.87 1.154 ;
      RECT 1.832 1.06 2.195 1.15 ;
      RECT 0.045 1.045 1.345 1.135 ;
      RECT 1.802 1.075 2.195 1.15 ;
      RECT 0.045 1.071 1.39 1.135 ;
  END
END AOI211X3H7R

MACRO AOI211X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211X4H7R 0 0 ;
  SIZE 3 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3 1.48 ;
        RECT 1.058 1.225 1.198 1.48 ;
        RECT 0.428 1.225 0.568 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3 0.08 ;
        RECT 2.478 -0.08 2.568 0.345 ;
        RECT 1.888 -0.08 2.028 0.185 ;
        RECT 1.233 -0.08 1.373 0.305 ;
        RECT 0.338 -0.08 0.428 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.348 0.855 1.248 0.945 ;
        RECT 1.158 0.637 1.248 0.945 ;
        RECT 0.348 0.638 0.438 0.945 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.693 0.655 0.993 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.023 0.455 2.175 0.655 ;
      LAYER MET2 ;
        RECT 2.05 0.23 2.15 0.76 ;
      LAYER VIA1 ;
        RECT 2.055 0.455 2.145 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.829 0.745 2.413 0.835 ;
        RECT 2.323 0.613 2.413 0.835 ;
        RECT 1.518 0.726 1.867 0.745 ;
        RECT 1.518 0.704 1.829 0.745 ;
        RECT 1.823 0.745 2.413 0.832 ;
        RECT 1.518 0.678 1.823 0.745 ;
        RECT 1.777 0.745 2.413 0.806 ;
        RECT 1.518 0.655 1.777 0.745 ;
        RECT 1.739 0.745 2.413 0.764 ;
        RECT 1.518 0.605 1.608 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.598 0.275 2.343 0.365 ;
        RECT 1.604 0.925 2.003 1.015 ;
        RECT 1.338 0.855 1.694 0.945 ;
        RECT 0.773 0.395 1.688 0.485 ;
        RECT 1.598 0.275 1.688 0.485 ;
        RECT 1.338 0.395 1.428 0.945 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.423 1.14 2.518 1.23 ;
      RECT 2.428 1.055 2.518 1.23 ;
      RECT 0.138 0.855 0.228 1.195 ;
      RECT 1.423 1.045 1.513 1.23 ;
      RECT 0.138 1.045 1.513 1.135 ;
  END
END AOI211X4H7R

MACRO AOI211X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211X6H7R 0 0 ;
  SIZE 4.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.6 1.48 ;
        RECT 1.9 1.225 2.04 1.48 ;
        RECT 1.37 1.225 1.51 1.48 ;
        RECT 0.84 1.225 0.98 1.48 ;
        RECT 0.31 1.225 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.6 0.08 ;
        RECT 4.3 -0.08 4.39 0.365 ;
        RECT 3.76 -0.08 3.9 0.185 ;
        RECT 3.23 -0.08 3.37 0.185 ;
        RECT 2.7 -0.08 2.84 0.185 ;
        RECT 2.14 -0.08 2.28 0.185 ;
        RECT 1.02 -0.08 1.16 0.185 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.02 0.51 2.11 0.65 ;
        RECT 0.2 0.51 2.11 0.6 ;
        RECT 0.2 0.455 0.375 0.6 ;
        RECT 0.2 0.455 0.29 0.65 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.74 1.865 0.83 ;
        RECT 0.425 0.74 0.575 0.945 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.45 0.69 4.265 0.78 ;
        RECT 2.38 0.655 2.575 0.733 ;
        RECT 2.38 0.526 2.47 0.733 ;
        RECT 2.426 0.69 4.265 0.768 ;
      LAYER MET2 ;
        RECT 2.45 0.6 2.55 1.135 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.76 0.51 3.975 0.6 ;
        RECT 3.825 0.455 3.975 0.6 ;
      LAYER MET2 ;
        RECT 3.85 0.23 3.95 0.76 ;
      LAYER VIA1 ;
        RECT 3.855 0.455 3.945 0.545 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.505 0.275 4.165 0.365 ;
        RECT 2.409 0.91 3.845 1 ;
        RECT 2.425 0.245 2.575 0.365 ;
        RECT 2.336 0.891 2.447 0.95 ;
        RECT 2.29 0.858 2.409 0.904 ;
        RECT 2.382 0.91 3.845 0.987 ;
        RECT 2.246 0.822 2.382 0.859 ;
        RECT 2.246 0.776 2.336 0.859 ;
        RECT 2.2 0.275 2.29 0.814 ;
      LAYER MET2 ;
        RECT 2.45 0.18 2.55 0.385 ;
      LAYER VIA1 ;
        RECT 2.455 0.255 2.545 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.328 1.09 4.34 1.18 ;
      RECT 4.25 1.035 4.34 1.18 ;
      RECT 2.321 1.048 2.328 1.177 ;
      RECT 2.283 1.09 4.34 1.154 ;
      RECT 0.045 1.045 2.321 1.135 ;
      RECT 0.045 1.071 2.366 1.135 ;
  END
END AOI211X6H7R

MACRO AOI21BX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21BX0P5H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.34 0.865 1.43 1.48 ;
        RECT 0.335 1.07 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.885 -0.08 0.975 0.415 ;
        RECT 0.07 -0.08 0.16 0.434 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.425 0.545 0.695 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.595 1.405 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.71 0.945 0.975 ;
        RECT 0.635 0.71 0.945 0.8 ;
        RECT 0.635 0.301 0.725 0.8 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.065 0.88 1.205 0.97 ;
      RECT 1.065 0.315 1.155 0.97 ;
      RECT 0.815 0.53 1.155 0.62 ;
      RECT 1.065 0.315 1.455 0.405 ;
      RECT 0.045 0.89 0.715 0.98 ;
  END
END AOI21BX0P5H7R

MACRO AOI21BX0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21BX0P7H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.34 0.897 1.43 1.48 ;
        RECT 0.335 1.07 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.885 -0.08 0.975 0.415 ;
        RECT 0.07 -0.08 0.16 0.425 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.425 0.545 0.695 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.595 1.405 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.71 0.945 0.975 ;
        RECT 0.635 0.71 0.945 0.8 ;
        RECT 0.635 0.3 0.725 0.8 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.065 0.85 1.205 0.94 ;
      RECT 1.065 0.334 1.155 0.94 ;
      RECT 0.815 0.53 1.155 0.62 ;
      RECT 1.065 0.334 1.44 0.424 ;
      RECT 0.045 0.89 0.715 0.98 ;
  END
END AOI21BX0P7H7R

MACRO AOI21BX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21BX1H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.34 0.945 1.43 1.48 ;
        RECT 0.335 1.07 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.885 -0.08 0.975 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.425 0.545 0.695 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.595 1.405 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.71 0.945 0.975 ;
        RECT 0.635 0.71 0.945 0.8 ;
        RECT 0.635 0.22 0.725 0.8 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.065 0.85 1.205 0.94 ;
      RECT 1.065 0.29 1.155 0.94 ;
      RECT 0.815 0.53 1.155 0.62 ;
      RECT 1.065 0.29 1.44 0.38 ;
      RECT 0.045 0.89 0.715 0.98 ;
  END
END AOI21BX1H7R

MACRO AOI21BX1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21BX1P4H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.34 0.989 1.43 1.48 ;
        RECT 0.335 1.07 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.885 -0.08 0.975 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.425 0.545 0.695 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.595 1.405 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.71 0.945 0.975 ;
        RECT 0.635 0.71 0.945 0.8 ;
        RECT 0.635 0.22 0.725 0.8 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.065 0.85 1.205 0.94 ;
      RECT 1.065 0.326 1.155 0.94 ;
      RECT 0.815 0.53 1.155 0.62 ;
      RECT 1.065 0.326 1.44 0.416 ;
      RECT 0.045 0.89 0.715 0.98 ;
  END
END AOI21BX1P4H7R

MACRO AOI21BX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21BX2H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.34 1.055 1.43 1.48 ;
        RECT 0.31 1.105 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.885 -0.08 0.975 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.425 0.545 0.695 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.625 1.435 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.745 0.945 0.975 ;
        RECT 0.635 0.745 0.945 0.835 ;
        RECT 0.635 0.22 0.725 0.835 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.065 0.85 1.205 0.94 ;
      RECT 1.065 0.36 1.155 0.94 ;
      RECT 0.815 0.565 1.155 0.655 ;
      RECT 1.065 0.36 1.315 0.45 ;
      RECT 0.045 0.925 0.715 1.015 ;
  END
END AOI21BX2H7R

MACRO AOI21BX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21BX3H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.555 1.015 1.695 1.48 ;
        RECT 0.31 1.115 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.555 -0.08 1.695 0.305 ;
        RECT 0.825 -0.08 0.965 0.305 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.425 0.545 0.695 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.51 0.655 1.81 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.635 0.395 1.19 0.485 ;
        RECT 1.1 0.28 1.19 0.485 ;
        RECT 0.85 0.755 0.945 0.975 ;
        RECT 0.635 0.755 0.945 0.845 ;
        RECT 0.635 0.245 0.725 0.845 ;
        RECT 0.575 0.245 0.725 0.335 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.83 0.835 1.92 0.98 ;
      RECT 1.33 0.28 1.42 0.98 ;
      RECT 1.33 0.835 1.92 0.925 ;
      RECT 0.895 0.575 1.42 0.665 ;
      RECT 1.33 0.395 1.92 0.485 ;
      RECT 1.83 0.28 1.92 0.485 ;
      RECT 0.625 1.065 1.19 1.155 ;
      RECT 1.1 0.96 1.19 1.155 ;
      RECT 0.625 0.935 0.715 1.155 ;
      RECT 0.045 0.935 0.715 1.025 ;
  END
END AOI21BX3H7R

MACRO AOI21BX4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21BX4H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.57 1.07 1.66 1.48 ;
        RECT 0.315 1.095 0.455 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.545 -0.08 1.685 0.305 ;
        RECT 0.815 -0.08 0.955 0.305 ;
        RECT 0.09 -0.08 0.18 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.57 0.545 0.795 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.5 0.655 1.8 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.635 0.395 1.18 0.485 ;
        RECT 1.09 0.345 1.18 0.485 ;
        RECT 0.814 0.855 0.975 0.945 ;
        RECT 0.725 0.836 0.852 0.879 ;
        RECT 0.725 0.795 0.814 0.879 ;
        RECT 0.771 0.855 0.975 0.924 ;
        RECT 0.681 0.751 0.771 0.834 ;
        RECT 0.635 0.345 0.725 0.789 ;
        RECT 0.565 0.345 0.725 0.435 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.32 0.875 1.935 0.965 ;
      RECT 1.32 0.355 1.41 0.965 ;
      RECT 0.885 0.575 1.41 0.665 ;
      RECT 1.32 0.395 1.91 0.485 ;
      RECT 1.82 0.318 1.91 0.485 ;
      RECT 0.545 1.065 1.205 1.155 ;
      RECT 0.545 0.91 0.635 1.155 ;
      RECT 0.09 0.91 0.18 1.05 ;
      RECT 0.09 0.91 0.635 1 ;
  END
END AOI21BX4H7R

MACRO AOI21BX6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21BX6H7R 0 0 ;
  SIZE 3 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3 1.48 ;
        RECT 2.552 1.055 2.642 1.48 ;
        RECT 2.052 1.07 2.142 1.48 ;
        RECT 0.547 1.095 0.687 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3 0.08 ;
        RECT 2.552 -0.08 2.642 0.345 ;
        RECT 2.027 -0.08 2.167 0.305 ;
        RECT 1.572 -0.08 1.662 0.345 ;
        RECT 1.047 -0.08 1.187 0.305 ;
        RECT 0.322 -0.08 0.412 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.625 0.475 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.65 0.58 0.785 0.78 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.982 0.655 2.522 0.745 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.987 0.855 1.687 0.945 ;
        RECT 0.797 0.395 1.437 0.485 ;
        RECT 0.987 0.395 1.077 0.945 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.802 0.875 2.417 0.965 ;
      RECT 1.802 0.355 1.892 0.965 ;
      RECT 1.167 0.625 1.892 0.715 ;
      RECT 1.802 0.395 2.417 0.485 ;
      RECT 0.797 1.065 1.437 1.155 ;
      RECT 0.797 0.915 0.887 1.155 ;
      RECT 0.297 0.915 0.887 1.005 ;
  END
END AOI21BX6H7R

MACRO AOI21X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X0P5H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.295 1.055 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.785 -0.08 0.925 0.175 ;
        RECT 0.07 -0.08 0.16 0.385 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.35 0.45 0.575 0.57 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.535 0.675 0.75 0.775 ;
        RECT 0.65 0.62 0.75 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.84 0.27 0.945 1.115 ;
        RECT 0.52 0.27 0.945 0.36 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.875 0.16 1.115 ;
      RECT 0.57 0.875 0.66 1.1 ;
      RECT 0.07 0.875 0.66 0.965 ;
  END
END AOI21X0P5H7R

MACRO AOI21X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X0P7H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.295 1.055 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.785 -0.08 0.925 0.185 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.35 0.455 0.575 0.575 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.52 0.68 0.75 0.775 ;
        RECT 0.655 0.625 0.75 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.84 0.275 0.945 1.083 ;
        RECT 0.52 0.275 0.945 0.365 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.875 0.16 1.083 ;
      RECT 0.57 0.875 0.66 1.068 ;
      RECT 0.07 0.875 0.66 0.965 ;
  END
END AOI21X0P7H7R

MACRO AOI21X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X1H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.31 1.055 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.785 -0.08 0.925 0.185 ;
        RECT 0.085 -0.08 0.175 0.385 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.455 0.575 0.545 ;
        RECT 0.425 0.455 0.525 0.68 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.64 0.625 0.76 0.775 ;
        RECT 0.67 0.525 0.76 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.97 0.945 1.11 ;
        RECT 0.855 0.275 0.945 1.11 ;
        RECT 0.52 0.275 0.945 0.365 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.085 0.87 0.175 1.035 ;
      RECT 0.585 0.87 0.675 1.02 ;
      RECT 0.085 0.87 0.675 0.96 ;
  END
END AOI21X1H7R

MACRO AOI21X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X1P4H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.785 -0.08 0.875 0.345 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.045 0.625 0.18 0.825 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 0.455 0.49 0.655 ;
        RECT 0.225 0.455 0.49 0.545 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.595 0.615 0.745 0.795 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.82 0.895 0.945 1.035 ;
        RECT 0.855 0.435 0.945 1.035 ;
        RECT 0.58 0.435 0.945 0.525 ;
        RECT 0.58 0.275 0.67 0.525 ;
        RECT 0.505 0.275 0.67 0.365 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.915 0.16 1.055 ;
      RECT 0.07 0.915 0.685 1.005 ;
  END
END AOI21X1P4H7R

MACRO AOI21X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X2H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.532 1.07 0.622 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.032 -0.08 1.172 0.185 ;
        RECT 0.282 -0.08 0.372 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.252 0.625 0.432 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.622 0.455 0.775 0.545 ;
        RECT 0.622 0.455 0.722 0.705 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.837 0.625 0.957 0.775 ;
        RECT 0.867 0.525 0.957 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.835 1.145 0.975 ;
        RECT 1.055 0.275 1.145 0.975 ;
        RECT 0.717 0.275 1.145 0.365 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.257 0.885 0.897 0.975 ;
  END
END AOI21X2H7R

MACRO AOI21X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X3H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.075 1.08 1.215 1.48 ;
        RECT 0.545 1.095 0.685 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.83 -0.08 1.92 0.345 ;
        RECT 1.33 -0.08 1.42 0.345 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.165 0.655 0.505 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.695 0.655 1.035 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.415 0.655 1.755 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.855 0.435 1.945 0.834 ;
        RECT 1.737 0.869 1.855 0.915 ;
        RECT 1.783 0.823 1.901 0.879 ;
        RECT 1.829 0.787 1.855 0.915 ;
        RECT 0.81 0.435 1.945 0.525 ;
        RECT 1.699 0.911 1.829 0.951 ;
        RECT 1.555 0.93 1.783 0.997 ;
        RECT 1.555 0.93 1.737 1.02 ;
        RECT 1.58 0.295 1.67 0.525 ;
        RECT 0.81 0.35 0.95 0.525 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.33 1.11 1.92 1.2 ;
      RECT 1.83 1.055 1.92 1.2 ;
      RECT 1.33 0.9 1.42 1.2 ;
      RECT 0.82 0.9 0.91 1.045 ;
      RECT 0.32 0.9 0.41 1.045 ;
      RECT 0.32 0.9 1.42 0.99 ;
      RECT 0.07 0.395 0.66 0.485 ;
      RECT 0.57 0.17 0.66 0.485 ;
      RECT 0.07 0.28 0.16 0.485 ;
      RECT 1.1 0.17 1.19 0.345 ;
      RECT 0.57 0.17 1.19 0.26 ;
  END
END AOI21X3H7R

MACRO AOI21X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X4H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 1.328 1.08 1.468 1.48 ;
        RECT 0.823 1.07 0.913 1.48 ;
        RECT 0.323 1.055 0.413 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 2.083 -0.08 2.173 0.345 ;
        RECT 1.583 -0.08 1.673 0.345 ;
        RECT 0.548 -0.08 0.688 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.418 0.655 0.758 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.948 0.655 1.288 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.625 0.655 1.965 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.055 0.435 2.145 0.887 ;
        RECT 1.808 0.885 2.101 0.932 ;
        RECT 1.997 0.866 2.145 0.887 ;
        RECT 2.035 0.837 2.055 0.965 ;
        RECT 1.063 0.435 2.145 0.525 ;
        RECT 1.808 0.885 2.035 0.975 ;
        RECT 1.833 0.37 1.923 0.525 ;
        RECT 1.063 0.395 1.203 0.525 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.583 1.065 2.198 1.155 ;
      RECT 1.583 0.885 1.673 1.155 ;
      RECT 0.548 0.885 1.673 0.975 ;
      RECT 0.323 0.395 0.913 0.485 ;
      RECT 0.823 0.205 0.913 0.485 ;
      RECT 0.323 0.28 0.413 0.485 ;
      RECT 1.353 0.205 1.443 0.345 ;
      RECT 0.823 0.205 1.443 0.295 ;
  END
END AOI21X4H7R

MACRO AOI21X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X6H7R 0 0 ;
  SIZE 3.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.2 1.48 ;
        RECT 1.787 1.08 1.927 1.48 ;
        RECT 1.282 1.07 1.372 1.48 ;
        RECT 0.782 1.07 0.872 1.48 ;
        RECT 0.282 1.055 0.372 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.2 0.08 ;
        RECT 2.542 -0.08 2.632 0.345 ;
        RECT 2.042 -0.08 2.132 0.345 ;
        RECT 0.757 -0.08 0.897 0.305 ;
        RECT 0.282 -0.08 0.372 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.427 0.655 0.967 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.182 0.655 1.722 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.162 0.655 2.702 0.745 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.267 0.875 2.882 0.965 ;
        RECT 2.792 0.286 2.882 0.965 ;
        RECT 1.257 0.455 2.882 0.545 ;
        RECT 2.292 0.37 2.382 0.545 ;
        RECT 1.787 0.38 1.927 0.545 ;
        RECT 1.257 0.395 1.397 0.545 ;
      LAYER MET2 ;
        RECT 2.05 0.23 2.15 0.76 ;
      LAYER VIA1 ;
        RECT 2.055 0.455 2.145 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.042 1.055 2.657 1.145 ;
      RECT 2.042 0.885 2.132 1.145 ;
      RECT 0.507 0.885 2.132 0.975 ;
      RECT 0.507 0.395 1.122 0.485 ;
      RECT 1.032 0.215 1.122 0.485 ;
      RECT 1.032 0.215 1.662 0.305 ;
  END
END AOI21X6H7R

MACRO AOI21X8H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X8H7R 0 0 ;
  SIZE 4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4 1.48 ;
        RECT 2.298 1.08 2.438 1.48 ;
        RECT 1.823 1.07 1.913 1.48 ;
        RECT 1.323 1.07 1.413 1.48 ;
        RECT 0.823 1.07 0.913 1.48 ;
        RECT 0.323 1.055 0.413 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4 0.08 ;
        RECT 3.553 -0.08 3.643 0.345 ;
        RECT 3.053 -0.08 3.143 0.33 ;
        RECT 2.553 -0.08 2.643 0.345 ;
        RECT 1.048 -0.08 1.188 0.305 ;
        RECT 0.548 -0.08 0.688 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.518 0.655 1.258 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.518 0.655 2.258 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.668 0.655 3.208 0.745 ;
      LAYER MET2 ;
        RECT 2.85 0.43 2.95 0.96 ;
      LAYER VIA1 ;
        RECT 2.855 0.655 2.945 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.778 0.865 3.393 0.955 ;
        RECT 3.303 0.37 3.393 0.955 ;
        RECT 2.098 0.455 3.393 0.545 ;
        RECT 2.803 0.37 2.893 0.545 ;
        RECT 1.548 0.395 2.188 0.485 ;
      LAYER MET2 ;
        RECT 2.65 0.23 2.75 0.76 ;
      LAYER VIA1 ;
        RECT 2.655 0.455 2.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.553 1.045 3.668 1.135 ;
      RECT 2.553 0.89 2.643 1.135 ;
      RECT 0.548 0.89 2.643 0.98 ;
      RECT 0.323 0.395 1.413 0.485 ;
      RECT 1.323 0.215 1.413 0.485 ;
      RECT 0.323 0.28 0.413 0.485 ;
      RECT 2.298 0.215 2.438 0.335 ;
      RECT 1.323 0.215 2.438 0.305 ;
  END
END AOI21X8H7R

MACRO AOI221X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221X0P5H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 0.335 1.14 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.535 -0.08 1.675 0.175 ;
        RECT 0.69 -0.08 0.83 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.6 0.59 0.8 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.31 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.625 1.035 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.195 0.455 1.375 0.545 ;
        RECT 1.195 0.455 1.285 0.665 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.445 0.625 1.545 0.895 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.64 0.275 1.745 1.06 ;
        RECT 0.095 0.275 1.745 0.365 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.805 1.14 1.475 1.23 ;
      RECT 0.045 0.96 1.21 1.05 ;
  END
END AOI221X0P5H7R

MACRO AOI221X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221X0P7H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 0.335 1.068 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.535 -0.08 1.675 0.175 ;
        RECT 0.69 -0.08 0.83 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.625 0.635 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.61 0.31 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.79 0.655 1.06 0.755 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.195 0.455 1.285 0.64 ;
        RECT 1.025 0.455 1.285 0.545 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.41 0.575 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.57 0.888 1.745 0.978 ;
        RECT 1.655 0.275 1.745 0.978 ;
        RECT 0.095 0.275 1.745 0.365 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.805 1.068 1.435 1.158 ;
      RECT 1.345 0.95 1.435 1.158 ;
      RECT 0.045 0.888 1.21 0.978 ;
  END
END AOI221X0P7H7R

MACRO AOI221X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221X1H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 0.335 1.14 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.535 -0.08 1.675 0.175 ;
        RECT 0.69 -0.08 0.83 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.575 0.59 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.605 0.31 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.605 1.035 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.195 0.455 1.375 0.545 ;
        RECT 1.195 0.455 1.285 0.665 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.445 0.605 1.545 0.875 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.64 0.275 1.745 1.06 ;
        RECT 0.095 0.275 1.745 0.365 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.805 1.14 1.475 1.23 ;
      RECT 0.045 0.96 1.21 1.05 ;
  END
END AOI221X1H7R

MACRO AOI221X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221X1P4H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 0.335 1.076 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.535 -0.08 1.675 0.175 ;
        RECT 0.69 -0.08 0.83 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.575 0.59 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.31 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.79 0.655 1.06 0.755 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.195 0.455 1.285 0.66 ;
        RECT 1.025 0.455 1.285 0.545 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.415 0.625 1.565 0.805 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.57 0.896 1.745 0.986 ;
        RECT 1.655 0.275 1.745 0.986 ;
        RECT 0.095 0.275 1.745 0.365 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.805 1.076 1.435 1.166 ;
      RECT 1.345 1.026 1.435 1.166 ;
      RECT 0.045 0.896 1.21 0.986 ;
  END
END AOI221X1P4H7R

MACRO AOI221X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221X2H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 0.537 1.07 0.627 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.787 -0.08 1.927 0.175 ;
        RECT 0.892 -0.08 1.032 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.64 0.6 0.82 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.615 0.512 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.625 1.265 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.397 0.455 1.59 0.545 ;
        RECT 1.397 0.455 1.487 0.715 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.655 0.615 1.76 0.885 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.85 0.275 1.96 0.975 ;
        RECT 0.297 0.275 1.96 0.365 ;
      LAYER MET2 ;
        RECT 1.85 0.625 1.95 1.16 ;
      LAYER VIA1 ;
        RECT 1.855 0.855 1.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.022 1.065 1.662 1.155 ;
      RECT 0.247 0.885 1.412 0.975 ;
  END
END AOI221X2H7R

MACRO AOI221X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221X3H7R 0 0 ;
  SIZE 3.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.2 1.48 ;
        RECT 1.045 1.095 1.185 1.48 ;
        RECT 0.545 1.095 0.685 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.2 0.08 ;
        RECT 2.6 -0.08 2.74 0.175 ;
        RECT 1.805 -0.08 1.945 0.175 ;
        RECT 1.06 -0.08 1.2 0.175 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.195 0.69 1.035 0.78 ;
        RECT 0.825 0.655 1.035 0.78 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.455 0.615 0.6 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.705 0.455 2.045 0.6 ;
      LAYER MET2 ;
        RECT 1.85 0.225 1.95 0.76 ;
      LAYER VIA1 ;
        RECT 1.855 0.455 1.945 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.44 0.69 2.295 0.78 ;
        RECT 2.205 0.636 2.295 0.78 ;
        RECT 1.225 0.655 1.515 0.745 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.565 0.63 2.855 0.77 ;
      LAYER MET2 ;
        RECT 2.65 0.43 2.75 0.96 ;
      LAYER VIA1 ;
        RECT 2.655 0.655 2.745 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.545 0.275 3.005 0.365 ;
        RECT 2.825 0.245 3.005 0.365 ;
        RECT 2.64 0.89 2.73 1.03 ;
        RECT 2.385 0.89 2.73 0.98 ;
        RECT 2.385 0.275 2.475 0.98 ;
      LAYER MET2 ;
        RECT 2.85 0.18 2.95 0.56 ;
      LAYER VIA1 ;
        RECT 2.855 0.255 2.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.29 1.14 2.98 1.23 ;
      RECT 2.89 1.035 2.98 1.23 ;
      RECT 0.82 0.905 0.91 1.045 ;
      RECT 0.32 0.905 0.41 1.045 ;
      RECT 0.32 0.905 2.225 1.005 ;
  END
END AOI221X3H7R

MACRO AOI221X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221X4H7R 0 0 ;
  SIZE 4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4 1.48 ;
        RECT 1.348 1.095 1.488 1.48 ;
        RECT 0.783 1.105 0.923 1.48 ;
        RECT 0.153 1.055 0.243 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4 0.08 ;
        RECT 3.203 -0.08 3.343 0.175 ;
        RECT 2.208 -0.08 2.348 0.175 ;
        RECT 1.363 -0.08 1.503 0.32 ;
        RECT 0.283 -0.08 0.373 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.231 0.64 1.375 0.745 ;
        RECT 0.333 0.745 1.254 0.757 ;
        RECT 1.126 0.726 1.375 0.745 ;
        RECT 1.21 0.65 1.231 0.779 ;
        RECT 0.333 0.745 1.21 0.812 ;
        RECT 1.164 0.684 1.375 0.745 ;
        RECT 0.333 0.745 1.164 0.835 ;
        RECT 0.333 0.64 0.423 0.835 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.565 0.988 0.655 ;
        RECT 0.625 0.455 0.775 0.655 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.155 0.565 2.498 0.655 ;
        RECT 2.225 0.455 2.375 0.655 ;
      LAYER MET2 ;
        RECT 2.25 0.23 2.35 0.76 ;
      LAYER VIA1 ;
        RECT 2.255 0.455 2.345 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.885 0.745 2.748 0.835 ;
        RECT 2.658 0.615 2.748 0.835 ;
        RECT 1.728 0.655 1.975 0.745 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.093 0.655 3.433 0.745 ;
      LAYER MET2 ;
        RECT 3.25 0.43 3.35 0.96 ;
      LAYER VIA1 ;
        RECT 3.255 0.655 3.345 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.643 0.275 3.658 0.365 ;
        RECT 2.855 0.885 3.308 0.975 ;
        RECT 2.855 0.275 2.945 0.975 ;
        RECT 1.112 0.41 1.733 0.5 ;
        RECT 1.643 0.275 1.733 0.5 ;
        RECT 1.112 0.275 1.202 0.5 ;
        RECT 0.848 0.275 1.202 0.365 ;
      LAYER MET2 ;
        RECT 2.85 0.23 2.95 0.76 ;
      LAYER VIA1 ;
        RECT 2.855 0.455 2.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.593 1.105 3.533 1.195 ;
      RECT 3.443 1.035 3.533 1.195 ;
      RECT 1.577 0.925 2.678 1.015 ;
      RECT 0.378 0.925 1.277 1.015 ;
      RECT 1.567 0.925 2.678 1.01 ;
      RECT 0.378 0.925 1.287 1.01 ;
      RECT 1.249 0.915 1.605 1.005 ;
      RECT 1.239 0.92 1.615 1.005 ;
  END
END AOI221X4H7R

MACRO AOI222X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222X0P5H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.29 -0.08 1.43 0.16 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.55 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.425 0.56 0.65 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.15 0.45 1.42 0.55 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.84 0.625 1.02 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.305 0.645 1.575 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.845 0.6 1.995 0.78 ;
      LAYER MET2 ;
        RECT 1.85 0.6 1.95 1.135 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.665 0.25 1.99 0.345 ;
        RECT 1.585 0.915 1.755 1.005 ;
        RECT 1.665 0.25 1.755 1.005 ;
        RECT 0.79 0.25 1.99 0.34 ;
      LAYER MET2 ;
        RECT 1.85 0.18 1.95 0.385 ;
      LAYER VIA1 ;
        RECT 1.855 0.255 1.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.57 0.915 0.66 1.155 ;
      RECT 0.07 0.915 0.16 1.155 ;
      RECT 0.07 0.915 1.195 1.005 ;
      RECT 0.79 1.095 1.99 1.185 ;
  END
END AOI222X0P5H7R

MACRO AOI222X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222X0P7H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.29 -0.08 1.43 0.16 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.55 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.425 0.56 0.65 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.185 0.455 1.375 0.545 ;
        RECT 1.185 0.455 1.275 0.655 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.84 0.625 1.02 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.44 0.615 1.575 0.815 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.845 0.6 1.995 0.78 ;
      LAYER MET2 ;
        RECT 1.85 0.6 1.95 1.135 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.665 0.25 1.99 0.345 ;
        RECT 1.585 0.915 1.755 1.005 ;
        RECT 1.665 0.25 1.755 1.005 ;
        RECT 0.79 0.25 1.99 0.34 ;
      LAYER MET2 ;
        RECT 1.85 0.18 1.95 0.385 ;
      LAYER VIA1 ;
        RECT 1.855 0.255 1.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.57 0.915 0.66 1.155 ;
      RECT 0.07 0.915 0.16 1.155 ;
      RECT 0.07 0.915 1.195 1.005 ;
      RECT 0.79 1.095 1.99 1.185 ;
  END
END AOI222X0P7H7R

MACRO AOI222X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222X1H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.29 -0.08 1.43 0.16 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.55 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.42 0.56 0.645 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.175 0.455 1.375 0.545 ;
        RECT 1.175 0.455 1.265 0.645 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.595 1.005 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.44 0.615 1.575 0.815 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.845 0.6 1.995 0.78 ;
      LAYER MET2 ;
        RECT 1.85 0.6 1.95 1.135 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.79 0.255 1.99 0.345 ;
        RECT 1.585 0.945 1.755 1.035 ;
        RECT 1.665 0.255 1.755 1.035 ;
      LAYER MET2 ;
        RECT 1.85 0.18 1.95 0.385 ;
      LAYER VIA1 ;
        RECT 1.855 0.255 1.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.79 1.14 1.99 1.23 ;
      RECT 1.85 1.095 1.99 1.23 ;
      RECT 1.32 1.095 1.46 1.23 ;
      RECT 0.79 1.095 0.93 1.23 ;
      RECT 0.57 0.915 0.66 1.075 ;
      RECT 0.07 0.915 0.16 1.075 ;
      RECT 1.055 0.915 1.195 1.035 ;
      RECT 0.07 0.915 1.195 1.005 ;
  END
END AOI222X1H7R

MACRO AOI222X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222X1P4H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.29 -0.08 1.43 0.305 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.55 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.425 0.555 0.695 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.175 0.595 1.345 0.785 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.595 1.005 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.595 1.585 0.815 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.855 0.6 2.015 0.78 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.625 0.255 2.02 0.345 ;
        RECT 1.605 0.905 1.765 0.995 ;
        RECT 1.675 0.255 1.765 0.995 ;
        RECT 1.04 0.415 1.765 0.505 ;
        RECT 1.625 0.255 1.765 0.505 ;
        RECT 1.04 0.255 1.13 0.505 ;
        RECT 0.79 0.255 1.13 0.345 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.56 ;
      LAYER VIA1 ;
        RECT 1.655 0.255 1.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.57 0.905 0.66 1.045 ;
      RECT 0.07 0.905 0.16 1.045 ;
      RECT 0.07 0.905 1.195 0.995 ;
      RECT 0.79 1.095 2.02 1.185 ;
  END
END AOI222X1P4H7R

MACRO AOI222X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222X2H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 0.533 1.07 0.623 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 1.553 -0.08 1.693 0.16 ;
        RECT 0.283 -0.08 0.373 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.55 0.545 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.425 0.755 0.705 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.388 0.455 1.575 0.545 ;
        RECT 1.388 0.455 1.478 0.68 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 0.595 1.2 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.625 0.64 1.883 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.158 0.625 2.345 0.775 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.803 0.255 2.303 0.345 ;
        RECT 1.898 0.835 2.063 0.925 ;
        RECT 1.973 0.255 2.063 0.925 ;
      LAYER MET2 ;
        RECT 1.85 0.18 1.95 0.56 ;
      LAYER VIA1 ;
        RECT 1.855 0.255 1.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.003 1.08 2.303 1.17 ;
      RECT 2.163 0.88 2.303 1.17 ;
      RECT 0.283 0.855 0.373 1.195 ;
      RECT 0.783 0.865 0.873 1.18 ;
      RECT 0.283 0.865 1.408 0.955 ;
  END
END AOI222X2H7R

MACRO AOI222X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222X3H7R 0 0 ;
  SIZE 3.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.6 1.48 ;
        RECT 1.045 1.095 1.185 1.48 ;
        RECT 0.545 1.095 0.685 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.6 0.08 ;
        RECT 2.885 -0.08 3.025 0.175 ;
        RECT 1.805 -0.08 1.945 0.175 ;
        RECT 1.06 -0.08 1.2 0.175 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.22 0.69 1.01 0.78 ;
        RECT 0.825 0.64 1.01 0.78 ;
        RECT 0.22 0.64 0.31 0.78 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.455 0.615 0.6 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.805 0.455 1.985 0.605 ;
      LAYER MET2 ;
        RECT 1.85 0.225 1.95 0.76 ;
      LAYER VIA1 ;
        RECT 1.855 0.455 1.945 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.695 2.295 0.785 ;
        RECT 2.205 0.64 2.295 0.785 ;
        RECT 1.455 0.625 1.545 0.785 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.8 0.455 2.98 0.605 ;
      LAYER MET2 ;
        RECT 2.85 0.23 2.95 0.76 ;
      LAYER VIA1 ;
        RECT 2.855 0.455 2.945 0.545 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.565 0.7 3.345 0.79 ;
        RECT 3.255 0.625 3.345 0.79 ;
        RECT 2.565 0.62 2.655 0.79 ;
      LAYER MET2 ;
        RECT 3.25 0.605 3.35 1.135 ;
      LAYER VIA1 ;
        RECT 3.255 0.655 3.345 0.745 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.545 0.275 3.525 0.365 ;
        RECT 3.225 0.255 3.375 0.365 ;
        RECT 3.145 0.895 3.235 1.04 ;
        RECT 2.385 0.895 3.235 0.985 ;
        RECT 2.64 0.895 2.73 1.04 ;
        RECT 2.385 0.275 2.475 0.985 ;
      LAYER MET2 ;
        RECT 3.25 0.18 3.35 0.385 ;
      LAYER VIA1 ;
        RECT 3.255 0.255 3.345 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.29 1.14 3.525 1.23 ;
      RECT 3.385 1.06 3.525 1.23 ;
      RECT 2.87 1.075 3.01 1.23 ;
      RECT 2.35 1.09 2.49 1.23 ;
      RECT 1.82 1.09 1.96 1.23 ;
      RECT 1.29 1.075 1.43 1.23 ;
      RECT 0.82 0.895 0.91 1.045 ;
      RECT 0.32 0.895 0.41 1.045 ;
      RECT 2.11 0.91 2.2 1.04 ;
      RECT 1.58 0.91 1.67 1.04 ;
      RECT 1.49 0.91 2.225 1 ;
      RECT 0.32 0.895 0.91 0.995 ;
      RECT 1.475 0.91 2.225 0.993 ;
      RECT 0.32 0.895 1.513 0.985 ;
      RECT 0.32 0.902 1.528 0.985 ;
  END
END AOI222X3H7R

MACRO AOI222X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222X4H7R 0 0 ;
  SIZE 4.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.6 1.48 ;
        RECT 1.453 1.11 1.593 1.48 ;
        RECT 0.823 1.11 0.963 1.48 ;
        RECT 0.283 1.055 0.373 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.6 0.08 ;
        RECT 3.578 -0.08 3.718 0.175 ;
        RECT 2.298 -0.08 2.438 0.175 ;
        RECT 1.453 -0.08 1.593 0.175 ;
        RECT 0.283 -0.08 0.373 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.433 0.745 1.345 0.835 ;
        RECT 1.255 0.615 1.345 0.835 ;
        RECT 0.433 0.615 0.523 0.835 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.688 0.565 1.028 0.655 ;
        RECT 0.825 0.455 0.975 0.655 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.225 0.565 2.565 0.655 ;
        RECT 2.225 0.455 2.375 0.655 ;
      LAYER MET2 ;
        RECT 2.25 0.23 2.35 0.76 ;
      LAYER VIA1 ;
        RECT 2.255 0.455 2.345 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.843 0.745 2.843 0.835 ;
        RECT 2.753 0.615 2.843 0.835 ;
        RECT 1.843 0.625 1.945 0.835 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.425 0.565 3.783 0.655 ;
        RECT 3.425 0.455 3.575 0.655 ;
      LAYER MET2 ;
        RECT 3.45 0.225 3.55 0.76 ;
      LAYER VIA1 ;
        RECT 3.455 0.455 3.545 0.545 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.153 0.745 4.145 0.835 ;
        RECT 4.055 0.615 4.145 0.835 ;
        RECT 3.153 0.615 3.243 0.835 ;
      LAYER MET2 ;
        RECT 4.05 0.43 4.15 0.96 ;
      LAYER VIA1 ;
        RECT 4.055 0.655 4.145 0.745 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.808 0.275 4.298 0.365 ;
        RECT 2.933 0.925 4.033 1.015 ;
        RECT 2.933 0.275 3.023 1.015 ;
        RECT 2.825 0.245 2.975 0.365 ;
      LAYER MET2 ;
        RECT 2.85 0.18 2.95 0.56 ;
      LAYER VIA1 ;
        RECT 2.855 0.255 2.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.683 1.11 4.273 1.2 ;
      RECT 4.183 1.055 4.273 1.2 ;
      RECT 0.503 0.925 2.768 1.015 ;
  END
END AOI222X4H7R

MACRO AOI22X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22X0P5H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.295 1.015 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.07 -0.08 1.16 0.355 ;
        RECT 0.045 -0.08 0.185 0.33 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.425 0.235 0.585 ;
      LAYER MET2 ;
        RECT 0.05 0.23 0.15 0.76 ;
      LAYER VIA1 ;
        RECT 0.055 0.455 0.145 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.312 0.655 0.612 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.425 0.76 0.575 ;
        RECT 0.565 0.425 0.76 0.55 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.55 1.155 0.82 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.795 0.945 0.945 1.035 ;
        RECT 0.855 0.225 0.945 1.035 ;
        RECT 0.545 0.225 0.945 0.315 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.56 ;
      LAYER VIA1 ;
        RECT 0.855 0.255 0.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.57 1.125 1.16 1.215 ;
      RECT 1.07 0.975 1.16 1.215 ;
      RECT 0.57 0.835 0.66 1.215 ;
      RECT 0.07 0.835 0.16 1.075 ;
      RECT 0.07 0.835 0.66 0.925 ;
  END
END AOI22X0P5H7R

MACRO AOI22X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22X0P7H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.295 1.045 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.07 -0.08 1.16 0.345 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.35 0.435 0.575 0.555 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 0.655 0.775 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.6 0.75 1.135 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.045 0.55 1.165 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.795 0.943 0.955 1.033 ;
        RECT 0.865 0.255 0.955 1.033 ;
        RECT 0.545 0.255 0.955 0.345 ;
      LAYER MET2 ;
        RECT 0.65 0.18 0.75 0.385 ;
      LAYER VIA1 ;
        RECT 0.655 0.255 0.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.57 1.123 1.16 1.213 ;
      RECT 1.07 1.005 1.16 1.213 ;
      RECT 0.57 0.865 0.66 1.213 ;
      RECT 0.07 0.865 0.16 1.073 ;
      RECT 0.07 0.865 0.66 0.955 ;
  END
END AOI22X0P7H7R

MACRO AOI22X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22X1H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.33 1.045 0.42 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.16 -0.08 1.25 0.345 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.43 0.39 0.55 0.615 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.165 0.625 1.345 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.64 0.625 0.82 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.91 0.255 1 1.035 ;
        RECT 0.635 0.255 1 0.345 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.56 ;
      LAYER VIA1 ;
        RECT 0.855 0.255 0.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.62 1.125 1.25 1.215 ;
      RECT 1.16 1.03 1.25 1.215 ;
      RECT 0.62 0.865 0.71 1.215 ;
      RECT 0.08 0.865 0.17 1.05 ;
      RECT 0.08 0.865 0.71 0.955 ;
  END
END AOI22X1H7R

MACRO AOI22X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22X1P4H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.33 1.045 0.42 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.16 -0.08 1.25 0.345 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.43 0.425 0.55 0.65 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.64 0.625 0.82 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.165 0.625 1.345 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.91 0.255 1 0.991 ;
        RECT 0.635 0.255 1 0.345 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.56 ;
      LAYER VIA1 ;
        RECT 0.855 0.255 0.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.62 1.081 1.25 1.171 ;
      RECT 1.16 1.03 1.25 1.171 ;
      RECT 0.62 0.865 0.71 1.171 ;
      RECT 0.08 0.865 0.17 1.006 ;
      RECT 0.08 0.865 0.71 0.955 ;
  END
END AOI22X1P4H7R

MACRO AOI22X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22X2H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 0.805 1.075 0.945 1.48 ;
        RECT 0.305 1.075 0.445 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 2.075 -0.08 2.215 0.345 ;
        RECT 1.085 -0.08 1.225 0.165 ;
        RECT 0.08 -0.08 0.17 0.37 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.495 0.655 1.835 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2 0.455 2.09 0.595 ;
        RECT 1.29 0.455 2.09 0.545 ;
        RECT 1.29 0.455 1.38 0.595 ;
      LAYER MET2 ;
        RECT 1.85 0.225 1.95 0.76 ;
      LAYER VIA1 ;
        RECT 1.855 0.455 1.945 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.93 0.455 1.02 0.6 ;
        RECT 0.23 0.455 1.02 0.545 ;
        RECT 0.23 0.455 0.32 0.6 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.655 0.795 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.23 0.895 2 0.985 ;
        RECT 0.555 0.255 1.74 0.345 ;
        RECT 1.23 0.715 1.32 0.985 ;
        RECT 1.11 0.715 1.32 0.805 ;
        RECT 1.11 0.255 1.2 0.805 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.56 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.035 1.075 2.265 1.165 ;
      RECT 0.07 0.895 0.16 1.135 ;
      RECT 0.58 0.895 0.67 1.12 ;
      RECT 1.035 0.895 1.125 1.165 ;
      RECT 0.07 0.895 1.125 0.985 ;
  END
END AOI22X2H7R

MACRO AOI22X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22X3H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 0.805 1.075 0.945 1.48 ;
        RECT 0.305 1.075 0.445 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 2.105 -0.08 2.245 0.345 ;
        RECT 1.085 -0.08 1.225 0.165 ;
        RECT 0.08 -0.08 0.17 0.37 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.03 0.455 2.12 0.655 ;
        RECT 1.29 0.455 2.12 0.545 ;
        RECT 1.29 0.455 1.38 0.63 ;
      LAYER MET2 ;
        RECT 1.85 0.225 1.95 0.76 ;
      LAYER VIA1 ;
        RECT 1.855 0.455 1.945 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.525 0.655 1.865 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.655 0.795 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.93 0.455 1.02 0.66 ;
        RECT 0.23 0.455 1.02 0.545 ;
        RECT 0.23 0.455 0.32 0.66 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.23 0.895 2.03 0.985 ;
        RECT 0.555 0.255 1.765 0.345 ;
        RECT 1.23 0.794 1.32 0.985 ;
        RECT 1.156 0.749 1.276 0.802 ;
        RECT 1.11 0.711 1.23 0.757 ;
        RECT 1.2 0.794 1.32 0.839 ;
        RECT 1.11 0.255 1.2 0.757 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.56 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.05 1.075 2.295 1.165 ;
      RECT 1.05 0.895 1.14 1.165 ;
      RECT 0.07 0.895 0.16 1.04 ;
      RECT 0.555 0.895 0.695 1.015 ;
      RECT 0.07 0.895 1.14 0.985 ;
  END
END AOI22X3H7R

MACRO AOI22X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22X4H7R 0 0 ;
  SIZE 4.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.6 1.48 ;
        RECT 1.91 1.225 2.05 1.48 ;
        RECT 1.38 1.225 1.52 1.48 ;
        RECT 0.85 1.225 0.99 1.48 ;
        RECT 0.32 1.225 0.46 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.6 0.08 ;
        RECT 4.33 -0.08 4.42 0.365 ;
        RECT 3.245 -0.08 3.385 0.175 ;
        RECT 2.195 -0.08 2.335 0.175 ;
        RECT 1.085 -0.08 1.225 0.175 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.65 0.655 3.805 0.745 ;
      LAYER MET2 ;
        RECT 2.85 0.43 2.95 0.96 ;
      LAYER VIA1 ;
        RECT 2.855 0.655 2.945 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.18 0.455 4.27 0.595 ;
        RECT 2.38 0.455 4.27 0.545 ;
        RECT 2.38 0.455 2.47 0.595 ;
      LAYER MET2 ;
        RECT 3.65 0.23 3.75 0.76 ;
      LAYER VIA1 ;
        RECT 3.655 0.455 3.745 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.485 0.655 1.845 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.02 0.455 2.11 0.595 ;
        RECT 0.235 0.455 2.11 0.545 ;
        RECT 0.235 0.455 0.325 0.595 ;
      LAYER MET2 ;
        RECT 1.65 0.23 1.75 0.76 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.2 0.855 4.18 0.955 ;
        RECT 0.555 0.265 3.875 0.355 ;
        RECT 2.2 0.265 2.29 0.955 ;
      LAYER MET2 ;
        RECT 4.05 0.63 4.15 1.16 ;
      LAYER VIA1 ;
        RECT 4.055 0.855 4.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 1.045 4.445 1.135 ;
  END
END AOI22X4H7R

MACRO AOI22X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22X6H7R 0 0 ;
  SIZE 4.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.6 1.48 ;
        RECT 1.91 1.225 2.05 1.48 ;
        RECT 1.38 1.1 1.52 1.48 ;
        RECT 0.85 1.1 0.99 1.48 ;
        RECT 0.32 1.1 0.46 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.6 0.08 ;
        RECT 4.305 -0.08 4.445 0.34 ;
        RECT 3.245 -0.08 3.385 0.175 ;
        RECT 2.195 -0.08 2.335 0.175 ;
        RECT 1.085 -0.08 1.225 0.175 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.865 0.69 3.985 0.78 ;
        RECT 2.615 0.655 2.955 0.745 ;
      LAYER MET2 ;
        RECT 2.65 0.43 2.75 0.96 ;
      LAYER VIA1 ;
        RECT 2.655 0.655 2.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.18 0.455 4.27 0.65 ;
        RECT 2.38 0.455 4.27 0.545 ;
        RECT 3.145 0.455 3.485 0.6 ;
        RECT 2.38 0.455 2.47 0.65 ;
      LAYER MET2 ;
        RECT 3.65 0.23 3.75 0.76 ;
      LAYER VIA1 ;
        RECT 3.655 0.455 3.745 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.735 0.69 1.845 0.78 ;
        RECT 0.485 0.655 0.825 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.02 0.455 2.11 0.65 ;
        RECT 0.23 0.455 2.11 0.545 ;
        RECT 0.985 0.455 1.325 0.6 ;
        RECT 0.23 0.455 0.32 0.65 ;
      LAYER MET2 ;
        RECT 1.65 0.23 1.75 0.76 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.2 0.895 4.18 0.985 ;
        RECT 0.585 0.265 3.875 0.355 ;
        RECT 2.2 0.825 2.345 0.985 ;
        RECT 2.2 0.265 2.29 0.985 ;
      LAYER MET2 ;
        RECT 2.25 0.63 2.35 1.16 ;
      LAYER VIA1 ;
        RECT 2.255 0.855 2.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.121 1.075 4.42 1.165 ;
      RECT 4.33 1.025 4.42 1.165 ;
      RECT 2.096 1.024 2.121 1.153 ;
      RECT 2.05 0.989 2.096 1.117 ;
      RECT 2.05 1.056 2.159 1.117 ;
      RECT 2.004 0.943 2.05 1.071 ;
      RECT 0.045 0.92 0.185 1.04 ;
      RECT 1.966 0.92 2.004 1.029 ;
      RECT 0.045 0.92 2.004 1.01 ;
  END
END AOI22X6H7R

MACRO AOI2BB1X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB1X0P5H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.575 1.215 0.715 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.12 -0.08 1.21 0.43 ;
        RECT 0.6 -0.08 0.69 0.355 ;
        RECT 0.07 -0.08 0.16 0.43 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.405 0.855 0.575 0.945 ;
        RECT 0.435 0.685 0.525 0.945 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.165 0.625 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 0.55 1.17 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.87 0.92 1.235 1.01 ;
        RECT 0.825 0.255 0.99 0.345 ;
        RECT 0.87 0.255 0.96 1.01 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.56 ;
      LAYER VIA1 ;
        RECT 0.855 0.255 0.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 1.035 0.775 1.125 ;
      RECT 0.685 0.445 0.775 1.125 ;
      RECT 0.07 0.935 0.16 1.125 ;
      RECT 0.32 0.445 0.775 0.535 ;
      RECT 0.32 0.305 0.41 0.535 ;
  END
END AOI2BB1X0P5H7R

MACRO AOI2BB1X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB1X0P7H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.575 1.215 0.715 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.12 -0.08 1.21 0.43 ;
        RECT 0.6 -0.08 0.69 0.355 ;
        RECT 0.07 -0.08 0.16 0.43 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.405 0.855 0.575 0.945 ;
        RECT 0.435 0.685 0.525 0.945 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.165 0.625 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 0.55 1.17 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.87 0.92 1.235 1.01 ;
        RECT 0.825 0.255 0.99 0.345 ;
        RECT 0.87 0.255 0.96 1.01 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.56 ;
      LAYER VIA1 ;
        RECT 0.855 0.255 0.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 1.035 0.775 1.125 ;
      RECT 0.685 0.445 0.775 1.125 ;
      RECT 0.07 0.935 0.16 1.125 ;
      RECT 0.32 0.445 0.775 0.535 ;
      RECT 0.32 0.305 0.41 0.535 ;
  END
END AOI2BB1X0P7H7R

MACRO AOI2BB1X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB1X1H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.575 1.215 0.715 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.12 -0.08 1.21 0.37 ;
        RECT 0.575 -0.08 0.715 0.345 ;
        RECT 0.07 -0.08 0.16 0.43 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.405 0.855 0.575 0.945 ;
        RECT 0.435 0.685 0.525 0.945 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.165 0.625 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 0.55 1.17 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.87 0.92 1.235 1.01 ;
        RECT 0.825 0.255 0.99 0.345 ;
        RECT 0.87 0.255 0.96 1.01 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.56 ;
      LAYER VIA1 ;
        RECT 0.855 0.255 0.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 1.035 0.775 1.125 ;
      RECT 0.685 0.445 0.775 1.125 ;
      RECT 0.07 0.935 0.16 1.125 ;
      RECT 0.32 0.445 0.775 0.535 ;
      RECT 0.32 0.305 0.41 0.535 ;
  END
END AOI2BB1X1H7R

MACRO AOI2BB1X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB1X1P4H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.575 1.215 0.715 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.12 -0.08 1.21 0.37 ;
        RECT 0.575 -0.08 0.715 0.345 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.405 0.855 0.575 0.945 ;
        RECT 0.435 0.66 0.525 0.945 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.165 0.625 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 0.55 1.17 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.87 0.92 1.235 1.01 ;
        RECT 0.825 0.255 0.99 0.345 ;
        RECT 0.87 0.255 0.96 1.01 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.56 ;
      LAYER VIA1 ;
        RECT 0.855 0.255 0.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 1.035 0.775 1.125 ;
      RECT 0.685 0.445 0.775 1.125 ;
      RECT 0.07 0.91 0.16 1.125 ;
      RECT 0.32 0.445 0.775 0.535 ;
      RECT 0.32 0.205 0.41 0.535 ;
  END
END AOI2BB1X1P4H7R

MACRO AOI2BB1X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB1X2H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.645 1.07 0.735 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.165 -0.08 1.255 0.345 ;
        RECT 0.645 -0.08 0.735 0.33 ;
        RECT 0.13 -0.08 0.22 0.345 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.755 0.575 0.98 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.36 0.825 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.095 0.655 1.395 0.745 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.165 0.855 1.255 1 ;
        RECT 0.915 0.855 1.255 0.945 ;
        RECT 0.915 0.37 1.005 0.945 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 1.04 0.245 1.13 ;
      RECT 0.045 0.445 0.135 1.13 ;
      RECT 0.73 0.445 0.82 0.705 ;
      RECT 0.045 0.445 0.82 0.535 ;
      RECT 0.38 0.22 0.47 0.535 ;
  END
END AOI2BB1X2H7R

MACRO AOI2BB1X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB1X3H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.08 1.06 1.22 1.48 ;
        RECT 0.56 1.225 0.7 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.605 -0.08 1.695 0.345 ;
        RECT 1.105 -0.08 1.195 0.33 ;
        RECT 0.585 -0.08 0.675 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.855 0.575 0.945 ;
        RECT 0.475 0.72 0.575 0.945 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.165 0.625 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.265 0.655 1.605 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.31 1.09 1.925 1.18 ;
        RECT 1.835 0.455 1.925 1.18 ;
        RECT 0.855 0.455 1.925 0.545 ;
        RECT 1.31 1.06 1.45 1.18 ;
        RECT 1.355 0.295 1.445 0.545 ;
        RECT 0.855 0.295 0.945 0.545 ;
      LAYER MET2 ;
        RECT 1.65 0.23 1.75 0.76 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.855 0.88 0.945 1.031 ;
      RECT 1.56 0.88 1.7 1 ;
      RECT 0.855 0.88 1.7 0.97 ;
      RECT 0.07 1.035 0.76 1.135 ;
      RECT 0.67 0.445 0.76 1.135 ;
      RECT 0.07 0.995 0.16 1.135 ;
      RECT 0.67 0.7 1.065 0.79 ;
      RECT 0.32 0.445 0.76 0.535 ;
      RECT 0.32 0.27 0.41 0.535 ;
  END
END AOI2BB1X3H7R

MACRO AOI2BB1X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB1X4H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.165 1.055 1.255 1.48 ;
        RECT 0.645 1.07 0.735 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.64 -0.08 1.78 0.305 ;
        RECT 1.14 -0.08 1.28 0.305 ;
        RECT 0.645 -0.08 0.735 0.33 ;
        RECT 0.13 -0.08 0.22 0.345 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.685 0.55 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.36 0.825 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.325 0.655 1.665 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.37 1.055 1.985 1.145 ;
        RECT 1.895 0.395 1.985 1.145 ;
        RECT 0.89 0.395 1.985 0.485 ;
      LAYER MET2 ;
        RECT 1.65 0.84 1.75 1.22 ;
      LAYER VIA1 ;
        RECT 1.655 1.055 1.745 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.92 0.245 1.01 ;
      RECT 0.045 0.445 0.135 1.01 ;
      RECT 0.685 0.625 1.1 0.715 ;
      RECT 0.685 0.445 0.775 0.715 ;
      RECT 0.045 0.445 0.775 0.535 ;
      RECT 0.38 0.32 0.47 0.535 ;
      RECT 0.89 0.865 1.76 0.955 ;
  END
END AOI2BB1X4H7R

MACRO AOI2BB1X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB1X6H7R 0 0 ;
  SIZE 2.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.8 1.48 ;
        RECT 1.327 1.07 1.417 1.48 ;
        RECT 0.822 1.07 0.912 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.8 0.08 ;
        RECT 2.302 -0.08 2.442 0.305 ;
        RECT 1.802 -0.08 1.942 0.305 ;
        RECT 1.302 -0.08 1.442 0.305 ;
        RECT 0.822 -0.08 0.912 0.33 ;
        RECT 0.322 -0.08 0.412 0.345 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.695 0.825 0.945 0.975 ;
        RECT 0.695 0.615 0.785 0.975 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.447 0.615 0.597 0.795 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.775 0.655 2.262 0.745 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.802 1.065 2.577 1.155 ;
        RECT 2.352 0.395 2.577 1.155 ;
        RECT 2.265 1.035 2.577 1.155 ;
        RECT 1.052 0.395 2.577 0.485 ;
      LAYER MET2 ;
        RECT 2.45 0.84 2.55 1.22 ;
      LAYER VIA1 ;
        RECT 2.455 1.055 2.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.267 0.885 0.437 0.975 ;
      RECT 0.267 0.435 0.357 0.975 ;
      RECT 1.016 0.625 1.407 0.715 ;
      RECT 1.002 0.58 1.016 0.708 ;
      RECT 0.956 0.55 1.002 0.678 ;
      RECT 0.91 0.504 0.956 0.632 ;
      RECT 0.91 0.606 1.054 0.632 ;
      RECT 0.864 0.458 0.91 0.586 ;
      RECT 0.826 0.504 0.956 0.544 ;
      RECT 0.267 0.435 0.864 0.525 ;
      RECT 0.572 0.37 0.662 0.525 ;
      RECT 1.052 0.885 2.192 0.975 ;
  END
END AOI2BB1X6H7R

MACRO AOI2BB2X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB2X0P5H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.29 1.16 1.38 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.485 -0.08 1.575 0.405 ;
        RECT 0.575 -0.08 0.715 0.185 ;
        RECT 0.07 -0.08 0.16 0.405 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.15 0.825 0.375 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.38 0.455 0.58 0.59 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.39 0.6 1.57 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.625 1.245 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.6 1.15 1.135 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.87 0.255 1.185 0.345 ;
        RECT 0.87 0.255 0.96 0.861 ;
        RECT 0.821 0.828 0.916 0.906 ;
        RECT 0.865 0.803 0.87 0.932 ;
        RECT 0.775 0.873 0.865 1.095 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.385 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.535 0.843 0.625 1.155 ;
      RECT 0.535 0.843 0.671 0.881 ;
      RECT 0.581 0.798 0.69 0.849 ;
      RECT 0.625 0.753 0.736 0.816 ;
      RECT 0.671 0.72 0.69 0.849 ;
      RECT 0.69 0.275 0.78 0.771 ;
      RECT 0.3 0.275 0.78 0.365 ;
      RECT 1 0.98 1.67 1.07 ;
  END
END AOI2BB2X0P5H7R

MACRO AOI2BB2X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB2X0P7H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.29 1.16 1.38 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.485 -0.08 1.575 0.405 ;
        RECT 0.575 -0.08 0.715 0.185 ;
        RECT 0.07 -0.08 0.16 0.405 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.15 0.825 0.375 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.38 0.455 0.58 0.59 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.39 0.625 1.57 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.625 1.245 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.6 1.15 1.135 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.87 0.255 1.175 0.345 ;
        RECT 0.87 0.255 0.96 0.861 ;
        RECT 0.821 0.828 0.916 0.906 ;
        RECT 0.865 0.803 0.87 0.932 ;
        RECT 0.775 0.873 0.865 1.095 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.385 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.535 0.843 0.625 1.155 ;
      RECT 0.535 0.843 0.671 0.881 ;
      RECT 0.581 0.798 0.69 0.849 ;
      RECT 0.625 0.753 0.736 0.816 ;
      RECT 0.671 0.72 0.69 0.849 ;
      RECT 0.69 0.275 0.78 0.771 ;
      RECT 0.3 0.275 0.78 0.365 ;
      RECT 1 0.98 1.67 1.07 ;
  END
END AOI2BB2X0P7H7R

MACRO AOI2BB2X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB2X1H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.29 1.16 1.38 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.485 -0.08 1.575 0.405 ;
        RECT 0.575 -0.08 0.715 0.185 ;
        RECT 0.07 -0.08 0.16 0.405 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.15 0.825 0.375 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.38 0.455 0.58 0.59 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.39 0.625 1.57 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.625 1.245 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.6 1.15 1.135 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.87 0.255 1.175 0.345 ;
        RECT 0.87 0.255 0.96 0.861 ;
        RECT 0.821 0.828 0.916 0.906 ;
        RECT 0.865 0.803 0.87 0.932 ;
        RECT 0.775 0.873 0.865 1.095 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.385 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.535 0.843 0.625 1.155 ;
      RECT 0.535 0.843 0.671 0.881 ;
      RECT 0.581 0.798 0.69 0.849 ;
      RECT 0.625 0.753 0.736 0.816 ;
      RECT 0.671 0.72 0.69 0.849 ;
      RECT 0.69 0.275 0.78 0.771 ;
      RECT 0.3 0.275 0.78 0.365 ;
      RECT 1 0.98 1.67 1.07 ;
  END
END AOI2BB2X1H7R

MACRO AOI2BB2X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB2X1P4H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.29 1.16 1.38 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.485 -0.08 1.575 0.405 ;
        RECT 0.575 -0.08 0.715 0.185 ;
        RECT 0.07 -0.08 0.16 0.405 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.15 0.825 0.375 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.38 0.455 0.58 0.59 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.375 0.625 1.57 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.625 1.245 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.6 1.15 1.135 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.87 0.255 1.175 0.345 ;
        RECT 0.87 0.255 0.96 0.861 ;
        RECT 0.821 0.828 0.916 0.906 ;
        RECT 0.865 0.803 0.87 0.932 ;
        RECT 0.775 0.873 0.865 1.095 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.385 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.535 0.843 0.625 1.155 ;
      RECT 0.535 0.843 0.671 0.881 ;
      RECT 0.581 0.798 0.69 0.849 ;
      RECT 0.625 0.753 0.736 0.816 ;
      RECT 0.671 0.72 0.69 0.849 ;
      RECT 0.69 0.275 0.78 0.771 ;
      RECT 0.3 0.275 0.78 0.365 ;
      RECT 1 0.98 1.67 1.07 ;
  END
END AOI2BB2X1P4H7R

MACRO AOI2BB2X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB2X2H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 2.13 1.225 2.27 1.48 ;
        RECT 1.6 1.225 1.74 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 2.44 -0.08 2.53 0.365 ;
        RECT 1.29 -0.08 1.38 0.35 ;
        RECT 0.705 -0.08 0.845 0.16 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.375 0.455 0.575 0.59 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.225 0.835 2.375 0.955 ;
        RECT 1.505 0.835 2.375 0.925 ;
      LAYER MET2 ;
        RECT 2.25 0.63 2.35 1.16 ;
      LAYER VIA1 ;
        RECT 2.255 0.855 2.345 0.945 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.765 0.655 2.105 0.745 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.01 0.455 1.98 0.545 ;
        RECT 1.89 0.24 1.98 0.545 ;
        RECT 1.04 0.865 1.415 0.955 ;
        RECT 1.325 0.455 1.415 0.955 ;
        RECT 1.01 0.24 1.1 0.545 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.57 0.825 0.66 1.155 ;
      RECT 0.57 0.825 0.755 0.915 ;
      RECT 0.665 0.265 0.755 0.915 ;
      RECT 0.665 0.635 1.235 0.725 ;
      RECT 0.295 0.265 0.755 0.355 ;
      RECT 0.775 1.045 2.545 1.135 ;
  END
END AOI2BB2X2H7R

MACRO AOI2BB2X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB2X3H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 2.13 1.225 2.27 1.48 ;
        RECT 1.6 1.225 1.74 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 2.42 -0.08 2.51 0.365 ;
        RECT 1.295 -0.08 1.385 0.35 ;
        RECT 0.705 -0.08 0.845 0.25 ;
        RECT 0.07 -0.08 0.16 0.39 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.365 0.625 0.545 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.485 0.7 2.385 0.79 ;
        RECT 2.225 0.655 2.385 0.79 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.795 0.51 2.135 0.6 ;
        RECT 1.795 0.455 1.975 0.6 ;
      LAYER MET2 ;
        RECT 1.85 0.225 1.95 0.76 ;
      LAYER VIA1 ;
        RECT 1.855 0.455 1.945 0.545 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.475 0.275 2.005 0.365 ;
        RECT 1.01 0.455 1.565 0.545 ;
        RECT 1.475 0.275 1.565 0.545 ;
        RECT 1.055 0.865 1.395 0.955 ;
        RECT 1.305 0.455 1.395 0.955 ;
        RECT 1.01 0.315 1.1 0.545 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.57 0.865 0.66 1.155 ;
      RECT 0.635 0.34 0.725 0.955 ;
      RECT 0.635 0.635 1.215 0.725 ;
      RECT 0.295 0.34 0.725 0.43 ;
      RECT 0.775 1.045 2.535 1.135 ;
  END
END AOI2BB2X3H7R

MACRO AOI2BB2X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB2X4H7R 0 0 ;
  SIZE 4.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.2 1.48 ;
        RECT 3.51 1.055 3.6 1.48 ;
        RECT 1.91 1.225 2.05 1.48 ;
        RECT 1.38 1.045 1.52 1.48 ;
        RECT 0.85 1.045 0.99 1.48 ;
        RECT 0.32 1.045 0.46 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.2 0.08 ;
        RECT 3.595 -0.08 3.735 0.305 ;
        RECT 2.72 -0.08 2.81 0.35 ;
        RECT 2.16 -0.08 2.3 0.175 ;
        RECT 1.085 -0.08 1.225 0.175 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.405 0.65 3.585 0.8 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.78 0.625 3.96 0.775 ;
      LAYER MET2 ;
        RECT 3.85 0.43 3.95 0.96 ;
      LAYER VIA1 ;
        RECT 3.855 0.655 3.945 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.03 0.455 2.12 0.595 ;
        RECT 0.23 0.455 2.12 0.545 ;
        RECT 0.23 0.455 0.32 0.595 ;
      LAYER MET2 ;
        RECT 1.65 0.23 1.75 0.76 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.49 0.655 1.875 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.255 0.895 3.11 0.985 ;
        RECT 0.585 0.265 2.585 0.355 ;
        RECT 2.255 0.265 2.345 0.985 ;
      LAYER MET2 ;
        RECT 2.25 0.63 2.35 1.16 ;
      LAYER VIA1 ;
        RECT 2.255 0.855 2.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 3.945 0.92 4.145 1.01 ;
      RECT 4.05 0.395 4.145 1.01 ;
      RECT 2.645 0.69 3.07 0.78 ;
      RECT 2.98 0.345 3.07 0.78 ;
      RECT 2.98 0.395 4.145 0.485 ;
      RECT 2.98 0.345 3.32 0.485 ;
      RECT 2.121 1.075 3.37 1.165 ;
      RECT 3.28 1.025 3.37 1.165 ;
      RECT 2.087 1.02 2.121 1.148 ;
      RECT 2.041 0.98 2.087 1.108 ;
      RECT 2.041 1.056 2.159 1.108 ;
      RECT 1.995 0.934 2.041 1.062 ;
      RECT 1.949 0.888 1.995 1.016 ;
      RECT 1.911 0.934 2.041 0.974 ;
      RECT 0.045 0.865 1.949 0.955 ;
  END
END AOI2BB2X4H7R

MACRO AOI2BB2X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB2X6H7R 0 0 ;
  SIZE 4.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.4 1.48 ;
        RECT 3.51 1.055 3.6 1.48 ;
        RECT 1.91 1.225 2.05 1.48 ;
        RECT 1.38 1.055 1.52 1.48 ;
        RECT 0.85 1.055 0.99 1.48 ;
        RECT 0.32 1.055 0.46 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.4 0.08 ;
        RECT 4.22 -0.08 4.31 0.365 ;
        RECT 3.695 -0.08 3.835 0.325 ;
        RECT 3.195 -0.08 3.335 0.325 ;
        RECT 2.68 -0.08 2.82 0.25 ;
        RECT 2.135 -0.08 2.275 0.175 ;
        RECT 1.085 -0.08 1.225 0.175 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.355 0.655 3.695 0.745 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.795 0.595 3.96 0.775 ;
      LAYER MET2 ;
        RECT 3.85 0.43 3.95 0.96 ;
      LAYER VIA1 ;
        RECT 3.855 0.655 3.945 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.02 0.455 2.11 0.65 ;
        RECT 0.23 0.455 2.11 0.545 ;
        RECT 0.985 0.455 1.325 0.6 ;
        RECT 0.23 0.455 0.32 0.65 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.75 0.69 1.845 0.78 ;
        RECT 0.485 0.655 0.825 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.2 0.895 3.11 0.985 ;
        RECT 2.2 0.34 3.085 0.43 ;
        RECT 2.2 0.855 2.375 0.985 ;
        RECT 2.2 0.265 2.29 0.985 ;
        RECT 0.555 0.265 2.29 0.355 ;
      LAYER MET2 ;
        RECT 2.25 0.63 2.35 1.16 ;
      LAYER VIA1 ;
        RECT 2.255 0.855 2.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 3.945 0.875 4.085 1.165 ;
      RECT 4.05 0.415 4.14 0.965 ;
      RECT 2.38 0.57 3.174 0.66 ;
      RECT 2.38 0.57 3.22 0.637 ;
      RECT 3.136 0.551 3.266 0.591 ;
      RECT 3.174 0.509 3.291 0.556 ;
      RECT 3.22 0.463 3.329 0.524 ;
      RECT 3.266 0.427 3.291 0.556 ;
      RECT 3.97 0.24 4.06 0.505 ;
      RECT 3.291 0.415 4.14 0.505 ;
      RECT 3.47 0.24 3.56 0.505 ;
      RECT 2.121 1.075 3.37 1.165 ;
      RECT 3.28 1.025 3.37 1.165 ;
      RECT 2.097 1.025 2.121 1.153 ;
      RECT 2.051 0.99 2.097 1.118 ;
      RECT 2.051 1.056 2.159 1.118 ;
      RECT 2.005 0.944 2.051 1.072 ;
      RECT 1.67 0.875 1.76 1.035 ;
      RECT 1.959 0.898 2.005 1.026 ;
      RECT 1.921 0.944 2.051 0.984 ;
      RECT 0.045 0.875 1.959 0.965 ;
  END
END AOI2BB2X6H7R

MACRO AOI2XB1X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2XB1X0P5H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.893 1.01 1.033 1.48 ;
        RECT 0.418 1.055 0.508 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.138 -0.08 1.278 0.175 ;
        RECT 0.418 -0.08 0.508 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.018 0.455 1.175 0.545 ;
        RECT 1.018 0.455 1.108 0.738 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END A0
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.44 0.45 0.56 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.588 1.365 0.823 ;
        RECT 1.265 0.525 1.365 0.823 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.403 0.96 1.545 1.05 ;
        RECT 1.455 0.27 1.545 1.05 ;
        RECT 0.643 0.27 1.545 0.36 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.168 0.932 1.258 1.095 ;
      RECT 0.648 0.83 0.738 1.075 ;
      RECT 1.134 0.847 1.168 0.975 ;
      RECT 1.096 0.887 1.214 0.939 ;
      RECT 0.648 0.83 1.134 0.92 ;
      RECT 0.045 1.04 0.283 1.13 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 0.045 0.65 0.883 0.74 ;
      RECT 0.045 0.23 0.283 0.32 ;
  END
END AOI2XB1X0P5H7R

MACRO AOI2XB1X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2XB1X0P7H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.893 1.042 1.033 1.48 ;
        RECT 0.418 1.055 0.508 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.138 -0.08 1.278 0.175 ;
        RECT 0.418 -0.08 0.508 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.018 0.455 1.175 0.545 ;
        RECT 1.018 0.455 1.108 0.721 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END A0
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.435 0.433 0.57 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.245 0.605 1.365 0.83 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.373 0.98 1.545 1.07 ;
        RECT 1.455 0.27 1.545 1.07 ;
        RECT 0.643 0.27 1.545 0.36 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.168 0.951 1.258 1.114 ;
      RECT 0.648 0.862 0.738 1.07 ;
      RECT 1.147 0.872 1.168 1.001 ;
      RECT 1.109 0.951 1.258 0.971 ;
      RECT 0.648 0.862 1.147 0.952 ;
      RECT 0.648 0.906 1.214 0.952 ;
      RECT 0.045 1.04 0.283 1.13 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 0.045 0.68 0.883 0.77 ;
      RECT 0.045 0.23 0.283 0.32 ;
  END
END AOI2XB1X0P7H7R

MACRO AOI2XB1X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2XB1X1H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.893 1.042 1.033 1.48 ;
        RECT 0.418 1.055 0.508 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.138 -0.08 1.278 0.175 ;
        RECT 0.418 -0.08 0.508 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.018 0.455 1.175 0.545 ;
        RECT 1.018 0.455 1.108 0.721 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END A0
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.435 0.433 0.57 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.245 0.605 1.365 0.83 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.373 0.98 1.545 1.07 ;
        RECT 1.455 0.27 1.545 1.07 ;
        RECT 0.643 0.27 1.545 0.36 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.168 0.951 1.258 1.114 ;
      RECT 0.648 0.862 0.738 1.07 ;
      RECT 1.147 0.872 1.168 1.001 ;
      RECT 1.109 0.951 1.258 0.971 ;
      RECT 0.648 0.862 1.147 0.952 ;
      RECT 0.648 0.906 1.214 0.952 ;
      RECT 0.045 1.04 0.283 1.13 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 0.045 0.68 0.883 0.77 ;
      RECT 0.045 0.23 0.283 0.32 ;
  END
END AOI2XB1X1H7R

MACRO AOI2XB1X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2XB1X1P4H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 0.892 1.095 1.032 1.48 ;
        RECT 0.418 1.055 0.508 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.168 -0.08 1.308 0.175 ;
        RECT 0.418 -0.08 0.508 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.455 1.175 0.545 ;
        RECT 1.025 0.455 1.118 0.73 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END A0
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.435 0.45 0.555 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.23 0.625 1.418 0.825 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.403 0.916 1.745 1.006 ;
        RECT 1.655 0.27 1.745 1.006 ;
        RECT 0.643 0.27 1.745 0.36 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.648 0.915 0.738 1.062 ;
      RECT 0.648 0.915 1.293 1.005 ;
      RECT 0.045 1.04 0.283 1.13 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 0.045 0.645 0.863 0.735 ;
      RECT 0.045 0.23 0.283 0.32 ;
  END
END AOI2XB1X1P4H7R

MACRO AOI2XB1X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2XB1X2H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 0.898 1.07 0.988 1.48 ;
        RECT 0.418 1.055 0.508 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.168 -0.08 1.308 0.175 ;
        RECT 0.393 -0.08 0.533 0.36 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.998 0.455 1.175 0.545 ;
        RECT 0.998 0.455 1.088 0.705 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END A0
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.45 0.45 0.57 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.225 0.625 1.425 0.76 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.425 0.85 1.623 0.945 ;
        RECT 1.533 0.27 1.623 0.945 ;
        RECT 0.643 0.27 1.623 0.36 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 1.04 0.283 1.13 ;
      RECT 0.045 0.27 0.135 1.13 ;
      RECT 0.045 0.66 0.838 0.75 ;
      RECT 0.748 0.61 0.838 0.75 ;
      RECT 0.045 0.27 0.283 0.36 ;
      RECT 0.623 0.865 1.263 0.955 ;
  END
END AOI2XB1X2H7R

MACRO AOI2XB1X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2XB1X3H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 1.623 1.095 1.763 1.48 ;
        RECT 1.123 1.095 1.263 1.48 ;
        RECT 0.648 1.055 0.738 1.48 ;
        RECT 0.418 1.055 0.508 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 2.158 -0.08 2.248 0.33 ;
        RECT 1.388 -0.08 1.528 0.175 ;
        RECT 0.418 -0.08 0.508 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.273 0.655 1.613 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A0
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.455 0.465 0.575 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.003 0.655 2.343 0.745 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.883 1.11 2.523 1.2 ;
        RECT 2.433 0.28 2.523 1.2 ;
        RECT 0.873 0.455 2.523 0.545 ;
        RECT 2.408 0.28 2.523 0.545 ;
        RECT 1.883 1.095 2.023 1.2 ;
        RECT 1.908 0.28 1.998 0.545 ;
        RECT 0.873 0.35 1.013 0.545 ;
      LAYER MET2 ;
        RECT 2.25 0.23 2.35 0.76 ;
      LAYER VIA1 ;
        RECT 2.255 0.455 2.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.898 0.915 0.988 1.055 ;
      RECT 1.373 0.915 1.513 1.035 ;
      RECT 2.133 0.915 2.273 1.02 ;
      RECT 0.898 0.915 2.273 1.005 ;
      RECT 0.648 0.17 0.738 0.375 ;
      RECT 1.123 0.265 1.793 0.355 ;
      RECT 1.123 0.17 1.213 0.355 ;
      RECT 0.648 0.17 1.213 0.26 ;
      RECT 0.045 0.98 0.283 1.07 ;
      RECT 0.045 0.23 0.135 1.07 ;
      RECT 0.045 0.665 1.063 0.755 ;
      RECT 0.045 0.23 0.283 0.32 ;
  END
END AOI2XB1X3H7R

MACRO AOI2XB1X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2XB1X4H7R 0 0 ;
  SIZE 3 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3 1.48 ;
        RECT 1.623 1.08 1.763 1.48 ;
        RECT 1.148 1.07 1.238 1.48 ;
        RECT 0.648 1.055 0.738 1.48 ;
        RECT 0.418 1.055 0.508 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3 0.08 ;
        RECT 2.258 -0.08 2.348 0.33 ;
        RECT 1.438 -0.08 1.578 0.175 ;
        RECT 0.418 -0.08 0.508 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.303 0.655 1.643 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A0
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.455 0.405 0.605 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.025 0.655 2.365 0.745 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.873 0.445 2.598 0.535 ;
        RECT 2.508 0.255 2.598 0.535 ;
        RECT 1.883 1.065 2.545 1.155 ;
        RECT 2.455 0.445 2.545 1.155 ;
        RECT 2.008 0.355 2.098 0.535 ;
        RECT 0.873 0.395 1.013 0.535 ;
      LAYER MET2 ;
        RECT 2.45 0.625 2.55 1.16 ;
      LAYER VIA1 ;
        RECT 2.455 0.855 2.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.148 0.265 1.893 0.355 ;
      RECT 0.648 0.215 0.738 0.355 ;
      RECT 0.648 0.215 1.238 0.305 ;
      RECT 0.045 0.92 0.283 1.01 ;
      RECT 0.045 0.275 0.135 1.01 ;
      RECT 0.045 0.695 0.571 0.785 ;
      RECT 0.045 0.695 0.611 0.764 ;
      RECT 0.573 0.655 1.063 0.745 ;
      RECT 0.533 0.676 1.063 0.745 ;
      RECT 0.571 0.656 0.573 0.784 ;
      RECT 0.045 0.275 0.283 0.365 ;
      RECT 0.873 0.885 2.273 0.975 ;
  END
END AOI2XB1X4H7R

MACRO AOI2XB1X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2XB1X6H7R 0 0 ;
  SIZE 3.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.6 1.48 ;
        RECT 1.997 1.095 2.137 1.48 ;
        RECT 1.487 1.095 1.627 1.48 ;
        RECT 0.987 1.095 1.127 1.48 ;
        RECT 0.532 1.055 0.622 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.6 0.08 ;
        RECT 2.892 -0.08 2.982 0.33 ;
        RECT 2.392 -0.08 2.482 0.33 ;
        RECT 1.802 -0.08 1.942 0.175 ;
        RECT 0.507 -0.08 0.647 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.597 0.655 2.337 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A0
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.425 0.545 0.695 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.51 0.655 3.05 0.745 ;
      LAYER MET2 ;
        RECT 2.65 0.43 2.75 0.96 ;
      LAYER VIA1 ;
        RECT 2.655 0.655 2.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.58 0.885 3.232 0.975 ;
        RECT 3.142 0.29 3.232 0.975 ;
        RECT 0.762 0.455 3.232 0.545 ;
        RECT 2.642 0.37 2.732 0.545 ;
        RECT 1.237 0.395 1.377 0.545 ;
        RECT 0.762 0.355 0.852 0.545 ;
      LAYER MET2 ;
        RECT 3.05 0.23 3.15 0.76 ;
      LAYER VIA1 ;
        RECT 3.055 0.455 3.145 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.297 1.065 2.97 1.155 ;
      RECT 2.297 0.915 2.387 1.155 ;
      RECT 0.737 0.915 2.387 1.005 ;
      RECT 1.537 0.265 2.257 0.355 ;
      RECT 0.987 0.215 1.627 0.305 ;
      RECT 0.257 0.85 0.56 0.94 ;
      RECT 0.257 0.85 0.606 0.917 ;
      RECT 0.522 0.831 0.652 0.871 ;
      RECT 0.257 0.245 0.347 0.94 ;
      RECT 0.56 0.789 0.652 0.871 ;
      RECT 0.56 0.789 0.698 0.825 ;
      RECT 0.606 0.743 0.717 0.793 ;
      RECT 0.606 0.743 0.755 0.764 ;
      RECT 0.717 0.655 1.377 0.745 ;
      RECT 0.652 0.697 1.377 0.745 ;
      RECT 0.698 0.664 0.717 0.793 ;
      RECT 0.257 0.245 0.397 0.335 ;
  END
END AOI2XB1X6H7R

MACRO AOI31X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31X0P5H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.58 0.76 0.725 0.985 ;
        RECT 0.1 0.76 0.725 0.85 ;
        RECT 0.1 0.76 0.19 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.155 -0.08 1.295 0.325 ;
        RECT 0.075 -0.08 0.215 0.325 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.425 0.235 0.58 ;
      LAYER MET2 ;
        RECT 0.05 0.23 0.15 0.76 ;
      LAYER VIA1 ;
        RECT 0.055 0.455 0.145 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.43 0.225 0.545 0.56 ;
      LAYER MET2 ;
        RECT 0.45 0.18 0.55 0.56 ;
      LAYER VIA1 ;
        RECT 0.455 0.255 0.545 0.345 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.425 0.835 0.575 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.165 0.425 1.345 0.58 ;
      LAYER MET2 ;
        RECT 1.25 0.18 1.35 0.585 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.12 0.77 1.345 0.985 ;
        RECT 0.975 0.77 1.345 0.86 ;
        RECT 0.975 0.225 1.065 0.86 ;
        RECT 0.845 0.225 1.065 0.315 ;
      LAYER MET2 ;
        RECT 1.25 0.815 1.35 1.22 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.325 1.105 0.975 1.195 ;
      RECT 0.835 0.95 0.975 1.195 ;
      RECT 0.325 0.94 0.465 1.195 ;
  END
END AOI31X0P5H7R

MACRO AOI31X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31X0P7H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.58 0.77 0.725 0.938 ;
        RECT 0.1 0.77 0.725 0.86 ;
        RECT 0.1 0.77 0.19 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.155 -0.08 1.295 0.325 ;
        RECT 0.075 -0.08 0.215 0.325 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.425 0.235 0.58 ;
      LAYER MET2 ;
        RECT 0.05 0.23 0.15 0.76 ;
      LAYER VIA1 ;
        RECT 0.055 0.455 0.145 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.225 0.545 0.585 ;
      LAYER MET2 ;
        RECT 0.45 0.18 0.55 0.56 ;
      LAYER VIA1 ;
        RECT 0.455 0.255 0.545 0.345 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.435 0.8 0.605 ;
        RECT 0.655 0.41 0.75 0.605 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.165 0.425 1.345 0.58 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.145 0.71 1.235 0.978 ;
        RECT 0.895 0.71 1.235 0.8 ;
        RECT 0.895 0.255 0.985 0.8 ;
        RECT 0.825 0.255 0.985 0.345 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.56 ;
      LAYER VIA1 ;
        RECT 0.855 0.255 0.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.325 1.03 0.95 1.12 ;
      RECT 0.86 0.925 0.95 1.12 ;
      RECT 0.325 0.95 0.465 1.12 ;
  END
END AOI31X0P7H7R

MACRO AOI31X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31X1H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.545 1.095 0.685 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.06 -0.08 1.2 0.35 ;
        RECT 0.07 -0.08 0.16 0.39 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.425 0.545 0.685 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.595 0.805 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.625 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.045 0.96 1.345 1.05 ;
        RECT 1.255 0.445 1.345 1.05 ;
        RECT 0.88 0.445 1.345 0.535 ;
        RECT 0.88 0.34 0.97 0.535 ;
        RECT 0.795 0.34 0.97 0.43 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.82 0.915 0.91 1.06 ;
      RECT 0.32 0.915 0.41 1.06 ;
      RECT 0.32 0.915 0.91 1.005 ;
  END
END AOI31X1H7R

MACRO AOI31X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31X1P4H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.545 1.095 0.685 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.135 -0.08 1.225 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.425 0.545 0.65 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.595 0.805 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.995 0.61 1.145 0.79 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.045 0.916 1.345 1.006 ;
        RECT 1.255 0.43 1.345 1.006 ;
        RECT 0.9 0.43 1.345 0.52 ;
        RECT 0.795 0.34 0.99 0.43 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.295 0.915 0.935 1.005 ;
  END
END AOI31X1P4H7R

MACRO AOI31X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31X2H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.755 1.07 0.845 1.48 ;
        RECT 0.255 1.055 0.345 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.19 -0.08 1.33 0.305 ;
        RECT 0.295 -0.08 0.385 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.625 0.445 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.635 0.425 0.745 0.705 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.595 1.005 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.165 0.625 1.345 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.23 0.885 1.545 0.975 ;
        RECT 1.455 0.395 1.545 0.975 ;
        RECT 0.94 0.395 1.545 0.485 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.48 0.89 1.12 0.98 ;
  END
END AOI31X2H7R

MACRO AOI31X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31X3H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 1.55 1.095 1.69 1.48 ;
        RECT 1.05 1.095 1.19 1.48 ;
        RECT 0.55 1.095 0.69 1.48 ;
        RECT 0.075 1.055 0.165 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 2.06 -0.08 2.2 0.335 ;
        RECT 0.3 -0.08 0.44 0.335 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.17 0.655 0.51 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.67 0.655 1.01 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.23 0.655 1.77 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.975 0.655 2.315 0.745 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.045 0.855 2.545 0.945 ;
        RECT 2.455 0.425 2.545 0.945 ;
        RECT 1.31 0.425 2.545 0.515 ;
        RECT 2.335 0.31 2.425 0.515 ;
        RECT 2.045 0.855 2.185 1.02 ;
        RECT 1.81 0.35 1.95 0.515 ;
        RECT 1.31 0.35 1.45 0.515 ;
      LAYER MET2 ;
        RECT 2.25 0.63 2.35 1.16 ;
      LAYER VIA1 ;
        RECT 2.255 0.855 2.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.82 1.11 2.41 1.2 ;
      RECT 2.32 1.055 2.41 1.2 ;
      RECT 1.82 0.915 1.91 1.2 ;
      RECT 1.3 0.915 1.44 1.035 ;
      RECT 0.8 0.915 0.94 1.035 ;
      RECT 0.3 0.915 0.44 1.035 ;
      RECT 0.3 0.915 1.91 1.005 ;
      RECT 1.56 0.17 1.7 0.335 ;
      RECT 0.8 0.17 0.94 0.335 ;
      RECT 0.8 0.17 1.7 0.26 ;
      RECT 0.07 0.425 1.19 0.515 ;
      RECT 1.05 0.35 1.19 0.515 ;
      RECT 0.575 0.325 0.665 0.515 ;
      RECT 0.07 0.31 0.16 0.515 ;
  END
END AOI31X3H7R

MACRO AOI31X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31X4H7R 0 0 ;
  SIZE 3 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3 1.48 ;
        RECT 1.757 1.095 1.897 1.48 ;
        RECT 1.257 1.095 1.397 1.48 ;
        RECT 0.757 1.095 0.897 1.48 ;
        RECT 0.272 1.055 0.362 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3 0.08 ;
        RECT 2.237 -0.08 2.377 0.305 ;
        RECT 0.507 -0.08 0.647 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.377 0.655 0.717 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.877 0.655 1.217 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.407 0.655 1.947 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.097 0.655 2.437 0.745 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.252 0.885 2.617 0.975 ;
        RECT 2.527 0.31 2.617 0.975 ;
        RECT 2.425 0.855 2.617 0.975 ;
        RECT 1.487 0.395 2.617 0.485 ;
        RECT 2.512 0.31 2.617 0.485 ;
        RECT 1.487 0.38 1.627 0.485 ;
      LAYER MET2 ;
        RECT 2.45 0.625 2.55 1.16 ;
      LAYER VIA1 ;
        RECT 2.455 0.855 2.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.027 1.08 2.642 1.17 ;
      RECT 2.027 0.915 2.117 1.17 ;
      RECT 0.507 0.915 2.117 1.005 ;
      RECT 1.737 0.2 1.877 0.305 ;
      RECT 1.007 0.2 1.147 0.305 ;
      RECT 1.007 0.2 1.877 0.29 ;
      RECT 0.277 0.395 1.397 0.485 ;
      RECT 1.257 0.38 1.397 0.485 ;
      RECT 0.277 0.31 0.367 0.485 ;
  END
END AOI31X4H7R

MACRO AOI32X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32X0P5H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.58 1.085 0.72 1.48 ;
        RECT 0.07 0.94 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.435 -0.08 1.525 0.345 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.43 0.425 0.55 0.65 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.645 0.595 0.795 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.435 0.62 1.555 0.845 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.065 0.455 1.375 0.545 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.15 0.91 1.29 1 ;
        RECT 1.15 0.655 1.24 1 ;
        RECT 0.885 0.655 1.24 0.745 ;
        RECT 0.885 0.245 0.975 0.745 ;
        RECT 0.835 0.245 0.975 0.335 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.91 1.09 1.525 1.18 ;
      RECT 1.435 0.94 1.525 1.18 ;
      RECT 0.91 0.905 1 1.18 ;
      RECT 0.32 0.905 0.41 1.045 ;
      RECT 0.32 0.905 1 0.995 ;
  END
END AOI32X0P5H7R

MACRO AOI32X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32X0P7H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.585 1.045 0.725 1.48 ;
        RECT 0.07 0.98 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.435 -0.08 1.525 0.345 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.43 0.425 0.55 0.65 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.595 0.805 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.435 0.59 1.555 0.815 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.095 0.425 1.345 0.58 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.15 0.958 1.29 1.048 ;
        RECT 1.15 0.67 1.24 1.048 ;
        RECT 0.895 0.67 1.24 0.76 ;
        RECT 0.895 0.255 0.985 0.76 ;
        RECT 0.825 0.255 0.985 0.345 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.56 ;
      LAYER VIA1 ;
        RECT 0.855 0.255 0.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.91 1.14 1.525 1.23 ;
      RECT 1.435 0.97 1.525 1.23 ;
      RECT 0.91 0.865 1 1.23 ;
      RECT 0.32 0.865 0.41 1.073 ;
      RECT 0.32 0.865 1 0.955 ;
  END
END AOI32X0P7H7R

MACRO AOI32X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32X1H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.545 1.095 0.685 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.36 -0.08 1.45 0.365 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.21 0.56 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.425 0.545 0.685 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.545 0.76 0.803 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.32 0.625 1.545 0.775 ;
        RECT 1.32 0.515 1.41 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.03 0.4 1.145 0.635 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.585 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.045 0.735 1.185 1.035 ;
        RECT 0.85 0.735 1.185 0.825 ;
        RECT 0.85 0.28 0.94 0.825 ;
        RECT 0.795 0.28 0.94 0.37 ;
      LAYER MET2 ;
        RECT 1.05 0.815 1.15 1.22 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.82 1.125 1.465 1.215 ;
      RECT 1.375 1.055 1.465 1.215 ;
      RECT 0.82 0.915 0.91 1.215 ;
      RECT 0.32 0.915 0.41 1.06 ;
      RECT 0.32 0.915 0.91 1.005 ;
  END
END AOI32X1H7R

MACRO AOI32X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32X1P4H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.545 1.095 0.685 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.36 -0.08 1.45 0.345 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.21 0.575 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.425 0.545 0.685 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.545 0.76 0.803 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.625 1.435 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.03 0.425 1.15 0.65 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.585 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.045 0.901 1.185 0.991 ;
        RECT 1.045 0.74 1.145 0.991 ;
        RECT 0.936 0.74 1.145 0.83 ;
        RECT 0.85 0.723 0.974 0.767 ;
        RECT 0.85 0.28 0.94 0.767 ;
        RECT 0.896 0.74 1.145 0.81 ;
        RECT 0.795 0.28 0.94 0.37 ;
      LAYER MET2 ;
        RECT 1.05 0.815 1.15 1.22 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.795 1.081 1.475 1.171 ;
      RECT 1.335 1.05 1.475 1.171 ;
      RECT 0.795 0.915 0.885 1.171 ;
      RECT 0.295 0.915 0.885 1.005 ;
  END
END AOI32X1P4H7R

MACRO AOI32X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32X2H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 0.757 1.095 0.897 1.48 ;
        RECT 0.282 1.055 0.372 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.572 -0.08 1.712 0.305 ;
        RECT 0.282 -0.08 0.372 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.575 0.545 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.425 0.745 0.725 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.6 0.99 0.8 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.505 0.645 1.775 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.125 0.645 1.395 0.745 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.257 0.855 1.955 0.945 ;
        RECT 1.865 0.395 1.955 0.945 ;
        RECT 1.007 0.395 1.955 0.485 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.032 1.035 1.712 1.125 ;
      RECT 1.032 0.915 1.122 1.125 ;
      RECT 0.507 0.915 1.122 1.005 ;
  END
END AOI32X2H7R

MACRO AOI32X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32X3H7R 0 0 ;
  SIZE 3.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.4 1.48 ;
        RECT 1.31 1.095 1.45 1.48 ;
        RECT 0.81 1.095 0.95 1.48 ;
        RECT 0.31 1.095 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.4 0.08 ;
        RECT 2.8 -0.08 2.94 0.335 ;
        RECT 0.295 -0.08 0.435 0.335 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.19 0.655 0.53 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.695 0.655 1.04 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.225 0.655 1.765 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.73 0.655 3.07 0.745 ;
      LAYER MET2 ;
        RECT 2.85 0.43 2.95 0.96 ;
      LAYER VIA1 ;
        RECT 2.855 0.655 2.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.925 0.655 2.265 0.745 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.8 0.855 2.94 1.02 ;
        RECT 2.055 0.855 2.94 0.945 ;
        RECT 2.36 0.35 2.45 0.945 ;
        RECT 1.305 0.425 2.45 0.515 ;
        RECT 2.305 0.35 2.45 0.515 ;
        RECT 2.055 0.855 2.195 1.02 ;
        RECT 1.805 0.35 1.945 0.515 ;
        RECT 1.305 0.35 1.445 0.515 ;
      LAYER MET2 ;
        RECT 2.45 0.625 2.55 1.16 ;
      LAYER VIA1 ;
        RECT 2.455 0.855 2.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.575 0.425 3.165 0.515 ;
      RECT 3.075 0.31 3.165 0.515 ;
      RECT 2.575 0.17 2.665 0.515 ;
      RECT 2.055 0.17 2.195 0.335 ;
      RECT 2.055 0.17 2.665 0.26 ;
      RECT 1.585 1.125 3.165 1.215 ;
      RECT 3.075 1.055 3.165 1.215 ;
      RECT 2.395 1.095 2.535 1.215 ;
      RECT 1.585 0.915 1.675 1.215 ;
      RECT 0.085 0.915 0.175 1.06 ;
      RECT 1.06 0.915 1.2 1.035 ;
      RECT 0.56 0.915 0.7 1.035 ;
      RECT 0.085 0.915 1.675 1.005 ;
      RECT 1.555 0.17 1.695 0.335 ;
      RECT 0.795 0.17 0.935 0.335 ;
      RECT 0.795 0.17 1.695 0.26 ;
      RECT 0.07 0.425 1.185 0.515 ;
      RECT 1.045 0.35 1.185 0.515 ;
      RECT 0.57 0.325 0.66 0.515 ;
      RECT 0.07 0.31 0.16 0.515 ;
  END
END AOI32X3H7R

MACRO AOI32X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32X4H7R 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.8 1.48 ;
        RECT 1.522 1.095 1.662 1.48 ;
        RECT 1.022 1.095 1.162 1.48 ;
        RECT 0.522 1.095 0.662 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.8 0.08 ;
        RECT 3.012 -0.08 3.152 0.305 ;
        RECT 0.507 -0.08 0.647 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.402 0.655 0.742 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.912 0.655 1.252 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.437 0.655 1.977 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.942 0.655 3.282 0.745 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.137 0.655 2.477 0.745 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.267 0.885 3.152 0.975 ;
        RECT 2.572 0.855 2.775 0.975 ;
        RECT 2.572 0.395 2.662 0.975 ;
        RECT 1.517 0.395 2.662 0.485 ;
      LAYER MET2 ;
        RECT 2.65 0.63 2.75 1.16 ;
      LAYER VIA1 ;
        RECT 2.655 0.855 2.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.797 1.065 3.402 1.155 ;
      RECT 1.797 0.915 1.887 1.155 ;
      RECT 0.272 0.915 1.887 1.005 ;
      RECT 2.787 0.395 3.377 0.485 ;
      RECT 3.287 0.31 3.377 0.485 ;
      RECT 2.787 0.215 2.877 0.485 ;
      RECT 2.267 0.215 2.877 0.305 ;
      RECT 0.282 0.395 1.397 0.485 ;
      RECT 0.282 0.31 0.372 0.485 ;
      RECT 1.007 0.215 1.907 0.305 ;
  END
END AOI32X4H7R

MACRO AOI33X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33X0P5H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 0.585 1.06 0.675 1.48 ;
        RECT 0.07 0.8 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.625 -0.08 1.715 0.335 ;
        RECT 0.045 -0.08 0.185 0.325 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.425 0.205 0.61 ;
      LAYER MET2 ;
        RECT 0.05 0.23 0.15 0.76 ;
      LAYER VIA1 ;
        RECT 0.055 0.455 0.145 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.415 0.4 0.545 0.61 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.49 0.75 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.505 0.425 1.745 0.585 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.585 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.225 1.36 0.61 ;
      LAYER MET2 ;
        RECT 1.25 0.18 1.35 0.56 ;
      LAYER VIA1 ;
        RECT 1.255 0.255 1.345 0.345 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.02 0.39 1.145 0.61 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.64 0.7 1.745 0.975 ;
        RECT 0.84 0.7 1.745 0.79 ;
        RECT 1.11 0.7 1.2 0.925 ;
        RECT 0.84 0.22 0.93 0.79 ;
      LAYER MET2 ;
        RECT 1.65 0.815 1.75 1.22 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.86 1.015 1.49 1.105 ;
      RECT 1.35 0.88 1.49 1.105 ;
      RECT 0.86 0.88 0.975 1.105 ;
      RECT 0.295 0.88 0.975 0.97 ;
  END
END AOI33X0P5H7R

MACRO AOI33X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33X0P7H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 0.585 1.045 0.675 1.48 ;
        RECT 0.07 0.89 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.61 -0.08 1.7 0.335 ;
        RECT 0.07 -0.08 0.16 0.35 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.41 0.545 0.61 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.505 0.755 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.565 0.425 1.745 0.575 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.585 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.225 1.345 0.585 ;
      LAYER MET2 ;
        RECT 1.25 0.18 1.35 0.56 ;
      LAYER VIA1 ;
        RECT 1.255 0.255 1.345 0.345 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.36 1.145 0.585 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.64 0.685 1.745 0.975 ;
        RECT 0.845 0.685 1.745 0.775 ;
        RECT 1.11 0.685 1.2 0.943 ;
        RECT 0.845 0.25 0.935 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.815 1.75 1.22 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.885 1.035 1.45 1.125 ;
      RECT 1.36 0.905 1.45 1.125 ;
      RECT 0.885 0.865 0.975 1.125 ;
      RECT 0.295 0.865 0.975 0.955 ;
  END
END AOI33X0P7H7R

MACRO AOI33X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33X1H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 0.585 1.135 0.675 1.48 ;
        RECT 0.07 0.925 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.59 -0.08 1.73 0.345 ;
        RECT 0.07 -0.08 0.16 0.4 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.62 0.255 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.435 0.425 0.545 0.671 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.505 0.755 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.54 1.64 0.63 ;
        RECT 1.455 0.425 1.545 0.63 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.225 1.35 0.655 ;
      LAYER MET2 ;
        RECT 1.25 0.18 1.35 0.56 ;
      LAYER VIA1 ;
        RECT 1.255 0.255 1.345 0.345 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.03 0.425 1.145 0.66 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.64 0.75 1.745 1 ;
        RECT 0.845 0.75 1.745 0.84 ;
        RECT 1.11 0.75 1.2 1.005 ;
        RECT 0.845 0.27 0.935 0.84 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.86 1.14 1.465 1.23 ;
      RECT 1.375 0.94 1.465 1.23 ;
      RECT 0.86 0.93 0.95 1.23 ;
      RECT 0.295 0.955 0.95 1.045 ;
  END
END AOI33X1H7R

MACRO AOI33X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33X1P4H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 0.585 1.1 0.675 1.48 ;
        RECT 0.07 0.969 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.615 -0.08 1.705 0.345 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.62 0.255 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.425 0.545 0.65 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.505 0.755 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.535 1.645 0.625 ;
        RECT 1.455 0.425 1.545 0.625 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.225 1.345 0.65 ;
      LAYER MET2 ;
        RECT 1.25 0.18 1.35 0.56 ;
      LAYER VIA1 ;
        RECT 1.255 0.255 1.345 0.345 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.425 1.145 0.65 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.64 0.74 1.745 1 ;
        RECT 0.845 0.74 1.745 0.83 ;
        RECT 1.085 0.74 1.225 0.905 ;
        RECT 0.845 0.315 0.935 0.83 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.86 0.995 1.475 1.085 ;
      RECT 0.295 0.92 0.95 1.01 ;
  END
END AOI33X1P4H7R

MACRO AOI33X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33X2H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 0.772 1.095 0.912 1.48 ;
        RECT 0.282 1.055 0.372 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.827 -0.08 1.917 0.345 ;
        RECT 0.282 -0.08 0.372 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.625 0.435 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.645 0.425 0.745 0.705 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.845 0.55 0.965 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.705 0.645 1.975 0.745 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.425 1.562 0.705 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.24 0.55 1.36 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.16 0.865 1.967 0.955 ;
        RECT 1.055 0.846 1.198 0.873 ;
        RECT 1.055 0.819 1.16 0.873 ;
        RECT 1.145 0.865 1.967 0.948 ;
        RECT 1.055 0.37 1.145 0.873 ;
        RECT 1.101 0.865 1.967 0.918 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.046 1.045 1.702 1.135 ;
      RECT 1.036 0.966 1.046 1.094 ;
      RECT 0.99 0.938 1.036 1.066 ;
      RECT 0.99 1.031 1.12 1.066 ;
      RECT 0.99 0.994 1.092 1.066 ;
      RECT 0.952 0.994 1.092 1.024 ;
      RECT 0.507 0.915 0.99 1.005 ;
  END
END AOI33X2H7R

MACRO AOI33X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33X3H7R 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.8 1.48 ;
        RECT 1.691 1.095 1.831 1.48 ;
        RECT 1.176 1.095 1.316 1.48 ;
        RECT 0.545 1.095 0.685 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.8 0.08 ;
        RECT 3.345 -0.08 3.485 0.335 ;
        RECT 0.295 -0.08 0.435 0.335 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.165 0.655 0.505 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.665 0.655 1.005 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.371 0.655 1.711 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.275 0.655 3.615 0.745 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.715 0.655 3.055 0.745 ;
      LAYER MET2 ;
        RECT 2.85 0.43 2.95 0.96 ;
      LAYER VIA1 ;
        RECT 2.855 0.655 2.945 0.745 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.955 0.655 2.295 0.745 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.345 0.855 3.485 1.02 ;
        RECT 2.186 0.855 3.485 0.945 ;
        RECT 2.845 0.855 2.985 1.02 ;
        RECT 2.385 0.35 2.475 0.945 ;
        RECT 1.305 0.44 2.475 0.53 ;
        RECT 2.335 0.35 2.475 0.53 ;
        RECT 2.186 0.855 2.326 1.02 ;
        RECT 1.82 0.32 1.96 0.53 ;
        RECT 1.305 0.35 1.445 0.53 ;
      LAYER MET2 ;
        RECT 2.465 0.63 2.565 1.16 ;
      LAYER VIA1 ;
        RECT 2.47 0.855 2.56 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.58 0.425 3.71 0.515 ;
      RECT 3.62 0.28 3.71 0.515 ;
      RECT 3.095 0.32 3.235 0.515 ;
      RECT 2.58 0.35 2.72 0.515 ;
      RECT 1.961 1.11 3.71 1.2 ;
      RECT 3.62 1.055 3.71 1.2 ;
      RECT 3.095 1.08 3.235 1.2 ;
      RECT 2.436 1.08 2.576 1.2 ;
      RECT 1.961 0.915 2.051 1.2 ;
      RECT 1.441 0.915 1.581 1.035 ;
      RECT 0.795 0.915 0.935 1.035 ;
      RECT 0.295 0.915 0.435 1.035 ;
      RECT 0.295 0.915 2.051 1.005 ;
      RECT 2.07 0.17 2.21 0.35 ;
      RECT 2.845 0.17 2.985 0.335 ;
      RECT 2.07 0.17 2.985 0.26 ;
      RECT 1.57 0.17 1.71 0.35 ;
      RECT 0.795 0.17 0.935 0.335 ;
      RECT 0.795 0.17 1.71 0.26 ;
      RECT 0.07 0.425 1.2 0.515 ;
      RECT 1.06 0.35 1.2 0.515 ;
      RECT 0.545 0.32 0.685 0.515 ;
      RECT 0.07 0.28 0.16 0.515 ;
  END
END AOI33X3H7R

MACRO AOI33X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33X4H7R 0 0 ;
  SIZE 4.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.2 1.48 ;
        RECT 1.888 1.095 2.028 1.48 ;
        RECT 1.388 1.095 1.528 1.48 ;
        RECT 0.757 1.095 0.897 1.48 ;
        RECT 0.282 1.055 0.372 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.2 0.08 ;
        RECT 3.527 -0.08 3.667 0.305 ;
        RECT 0.507 -0.08 0.647 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.377 0.655 0.717 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.877 0.655 1.217 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.568 0.655 1.908 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.457 0.655 3.797 0.745 ;
      LAYER MET2 ;
        RECT 3.65 0.43 3.75 0.96 ;
      LAYER VIA1 ;
        RECT 3.655 0.655 3.745 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.897 0.655 3.237 0.745 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.152 0.655 2.492 0.745 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.383 0.885 3.667 0.975 ;
        RECT 2.655 0.575 2.745 0.975 ;
        RECT 2.582 0.38 2.672 0.665 ;
        RECT 1.502 0.395 2.672 0.485 ;
        RECT 2.532 0.38 2.672 0.485 ;
        RECT 1.502 0.38 1.642 0.485 ;
      LAYER MET2 ;
        RECT 2.65 0.43 2.75 0.96 ;
      LAYER VIA1 ;
        RECT 2.655 0.655 2.745 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.158 1.065 3.917 1.155 ;
      RECT 2.158 0.915 2.248 1.155 ;
      RECT 0.507 0.915 2.248 1.005 ;
      RECT 2.762 0.395 3.892 0.485 ;
      RECT 3.802 0.28 3.892 0.485 ;
      RECT 2.762 0.38 2.902 0.485 ;
      RECT 3.027 0.2 3.167 0.305 ;
      RECT 2.267 0.2 2.407 0.305 ;
      RECT 2.267 0.2 3.167 0.29 ;
      RECT 1.767 0.2 1.907 0.305 ;
      RECT 1.007 0.2 1.147 0.305 ;
      RECT 1.007 0.2 1.907 0.29 ;
      RECT 0.282 0.395 1.412 0.485 ;
      RECT 1.272 0.38 1.412 0.485 ;
      RECT 0.282 0.28 0.372 0.485 ;
  END
END AOI33X4H7R

MACRO BUFX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX0P5H7R 0 0 ;
  SIZE 0.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.8 1.48 ;
        RECT 0.325 1.07 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.8 0.08 ;
        RECT 0.325 -0.08 0.415 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.43 0.575 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.555 1.065 0.745 1.155 ;
        RECT 0.655 0.23 0.745 1.155 ;
        RECT 0.555 0.23 0.745 0.32 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.205 0.16 1.155 ;
      RECT 0.07 0.79 0.545 0.88 ;
  END
END BUFX0P5H7R

MACRO BUFX0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX0P7H7R 0 0 ;
  SIZE 0.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.8 1.48 ;
        RECT 0.325 1.07 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.8 0.08 ;
        RECT 0.325 -0.08 0.415 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.755 0.375 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.58 0.225 0.745 0.375 ;
        RECT 0.58 0.225 0.67 1.123 ;
      LAYER MET2 ;
        RECT 0.65 0.18 0.75 0.56 ;
      LAYER VIA1 ;
        RECT 0.655 0.255 0.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.205 0.16 1.155 ;
      RECT 0.07 0.465 0.49 0.605 ;
  END
END BUFX0P7H7R

MACRO BUFX10H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX10H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 1.82 1.07 1.91 1.48 ;
        RECT 1.32 1.07 1.41 1.48 ;
        RECT 0.82 1.07 0.91 1.48 ;
        RECT 0.32 1.055 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 2.32 -0.08 2.41 0.345 ;
        RECT 1.795 -0.08 1.935 0.305 ;
        RECT 1.295 -0.08 1.435 0.305 ;
        RECT 0.795 -0.08 0.935 0.305 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.655 0.765 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.07 0.22 2.16 1.165 ;
        RECT 1.07 0.855 2.16 0.945 ;
        RECT 1.045 0.395 2.16 0.485 ;
        RECT 1.57 0.855 1.66 1.17 ;
        RECT 1.07 0.855 1.16 1.21 ;
      LAYER MET2 ;
        RECT 1.85 0.625 1.95 1.16 ;
      LAYER VIA1 ;
        RECT 1.855 0.855 1.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.545 0.885 0.945 0.975 ;
      RECT 0.855 0.395 0.945 0.975 ;
      RECT 0.855 0.625 1.915 0.715 ;
      RECT 0.07 0.395 0.945 0.485 ;
      RECT 0.57 0.27 0.66 0.485 ;
      RECT 0.07 0.255 0.16 0.485 ;
  END
END BUFX10H7R

MACRO BUFX12H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX12H7R 0 0 ;
  SIZE 2.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.8 1.48 ;
        RECT 2.32 1.055 2.41 1.48 ;
        RECT 1.82 1.07 1.91 1.48 ;
        RECT 1.32 1.07 1.41 1.48 ;
        RECT 0.82 1.07 0.91 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.8 0.08 ;
        RECT 2.295 -0.08 2.435 0.305 ;
        RECT 1.795 -0.08 1.935 0.305 ;
        RECT 1.295 -0.08 1.435 0.305 ;
        RECT 0.795 -0.08 0.935 0.305 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.655 0.765 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.07 0.855 2.66 0.945 ;
        RECT 2.57 0.205 2.66 0.945 ;
        RECT 1.045 0.395 2.66 0.485 ;
        RECT 2.07 0.855 2.16 1.17 ;
        RECT 2.07 0.22 2.16 0.485 ;
        RECT 1.57 0.855 1.66 1.17 ;
        RECT 1.07 0.855 1.16 1.21 ;
      LAYER MET2 ;
        RECT 2.45 0.625 2.55 1.16 ;
      LAYER VIA1 ;
        RECT 2.455 0.855 2.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.885 0.16 1.175 ;
      RECT 0.07 0.885 0.945 0.975 ;
      RECT 0.855 0.395 0.945 0.975 ;
      RECT 0.855 0.625 2.315 0.715 ;
      RECT 0.07 0.395 0.945 0.485 ;
      RECT 0.07 0.205 0.16 0.485 ;
  END
END BUFX12H7R

MACRO BUFX16H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX16H7R 0 0 ;
  SIZE 3.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.6 1.48 ;
        RECT 3.075 0.855 3.165 1.48 ;
        RECT 2.575 1.07 2.665 1.48 ;
        RECT 2.075 1.07 2.165 1.48 ;
        RECT 1.575 1.07 1.665 1.48 ;
        RECT 1.075 1.07 1.165 1.48 ;
        RECT 0.575 1.07 0.665 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.6 0.08 ;
        RECT 3.075 -0.08 3.165 0.345 ;
        RECT 2.55 -0.08 2.69 0.305 ;
        RECT 2.05 -0.08 2.19 0.305 ;
        RECT 1.55 -0.08 1.69 0.305 ;
        RECT 1.05 -0.08 1.19 0.305 ;
        RECT 0.55 -0.08 0.69 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.47 0.655 1.01 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.825 0.395 2.94 1.15 ;
        RECT 1.325 0.855 2.94 0.945 ;
        RECT 1.3 0.395 2.94 0.485 ;
        RECT 2.325 0.855 2.415 1.17 ;
        RECT 1.825 0.855 1.915 1.17 ;
        RECT 1.325 0.855 1.415 1.21 ;
      LAYER MET2 ;
        RECT 2.65 0.63 2.75 1.16 ;
      LAYER VIA1 ;
        RECT 2.655 0.855 2.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.825 0.855 0.915 1.005 ;
      RECT 0.3 0.855 1.19 0.945 ;
      RECT 1.1 0.395 1.19 0.945 ;
      RECT 1.1 0.625 2.57 0.715 ;
      RECT 0.325 0.395 1.19 0.485 ;
      RECT 0.325 0.345 0.415 0.485 ;
  END
END BUFX16H7R

MACRO BUFX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX1H7R 0 0 ;
  SIZE 0.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.8 1.48 ;
        RECT 0.325 1.07 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.8 0.08 ;
        RECT 0.325 -0.08 0.415 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.745 0.37 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.555 1.045 0.745 1.135 ;
        RECT 0.655 0.265 0.745 1.135 ;
        RECT 0.555 0.265 0.745 0.355 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.205 0.16 1.155 ;
      RECT 0.07 0.5 0.545 0.59 ;
  END
END BUFX1H7R

MACRO BUFX1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX1P4H7R 0 0 ;
  SIZE 0.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.8 1.48 ;
        RECT 0.325 1.07 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.8 0.08 ;
        RECT 0.325 -0.08 0.415 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.58 0.825 0.745 1.031 ;
        RECT 0.58 0.301 0.67 1.031 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.865 0.16 1.155 ;
      RECT 0.07 0.865 0.49 0.955 ;
      RECT 0.4 0.435 0.49 0.955 ;
      RECT 0.07 0.435 0.49 0.525 ;
      RECT 0.07 0.205 0.16 0.525 ;
  END
END BUFX1P4H7R

MACRO BUFX20H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX20H7R 0 0 ;
  SIZE 4.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.4 1.48 ;
        RECT 3.825 0.855 3.915 1.48 ;
        RECT 3.325 1.07 3.415 1.48 ;
        RECT 2.825 1.07 2.915 1.48 ;
        RECT 2.325 1.07 2.415 1.48 ;
        RECT 1.825 1.07 1.915 1.48 ;
        RECT 1.325 1.07 1.415 1.48 ;
        RECT 0.825 1.07 0.915 1.48 ;
        RECT 0.325 0.855 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.4 0.08 ;
        RECT 3.8 -0.08 3.94 0.305 ;
        RECT 3.3 -0.08 3.44 0.305 ;
        RECT 2.8 -0.08 2.94 0.305 ;
        RECT 2.3 -0.08 2.44 0.305 ;
        RECT 1.8 -0.08 1.94 0.305 ;
        RECT 1.3 -0.08 1.44 0.305 ;
        RECT 0.8 -0.08 0.94 0.305 ;
        RECT 0.325 -0.08 0.415 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.48 0.655 1.22 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.55 0.395 4.165 0.485 ;
        RECT 4.075 0.255 4.165 0.485 ;
        RECT 3.575 0.395 3.665 1.165 ;
        RECT 1.575 0.855 3.665 0.945 ;
        RECT 3.075 0.855 3.165 1.17 ;
        RECT 2.575 0.855 2.665 1.17 ;
        RECT 2.075 0.855 2.165 1.17 ;
        RECT 1.575 0.855 1.665 1.21 ;
      LAYER MET2 ;
        RECT 3.45 0.625 3.55 1.16 ;
      LAYER VIA1 ;
        RECT 3.455 0.855 3.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.885 1.4 0.975 ;
      RECT 1.31 0.395 1.4 0.975 ;
      RECT 1.31 0.625 3.42 0.715 ;
      RECT 0.55 0.395 1.4 0.485 ;
  END
END BUFX20H7R

MACRO BUFX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX2H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.325 1.07 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.325 -0.08 0.415 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.165 0.625 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.555 1.045 0.745 1.135 ;
        RECT 0.655 0.265 0.745 1.135 ;
        RECT 0.555 0.265 0.745 0.355 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.865 0.16 1.155 ;
      RECT 0.07 0.865 0.565 0.955 ;
      RECT 0.475 0.445 0.565 0.955 ;
      RECT 0.07 0.445 0.565 0.535 ;
      RECT 0.07 0.205 0.16 0.535 ;
  END
END BUFX2H7R

MACRO BUFX2P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX2P5H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.835 1.055 0.925 1.48 ;
        RECT 0.325 1.07 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.835 -0.08 0.925 0.345 ;
        RECT 0.325 -0.08 0.415 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.555 1.065 0.745 1.155 ;
        RECT 0.655 0.23 0.745 1.155 ;
        RECT 0.555 0.23 0.745 0.32 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.865 0.16 1.155 ;
      RECT 0.07 0.865 0.565 0.955 ;
      RECT 0.475 0.435 0.565 0.955 ;
      RECT 0.07 0.435 0.565 0.525 ;
      RECT 0.07 0.205 0.16 0.525 ;
  END
END BUFX2P5H7R

MACRO BUFX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX3H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.835 1.055 0.925 1.48 ;
        RECT 0.325 1.07 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.835 -0.08 0.925 0.345 ;
        RECT 0.325 -0.08 0.415 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.165 0.625 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.555 1.045 0.745 1.135 ;
        RECT 0.655 0.245 0.745 1.135 ;
        RECT 0.555 0.245 0.745 0.335 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.865 0.16 1.155 ;
      RECT 0.07 0.865 0.549 0.955 ;
      RECT 0.459 0.445 0.549 0.955 ;
      RECT 0.07 0.445 0.549 0.535 ;
      RECT 0.07 0.205 0.16 0.535 ;
  END
END BUFX3H7R

MACRO BUFX3P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX3P5H7R 0 0 ;
  SIZE 1.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.2 1.48 ;
        RECT 0.835 1.055 0.925 1.48 ;
        RECT 0.325 1.07 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.2 0.08 ;
        RECT 0.835 -0.08 0.925 0.345 ;
        RECT 0.325 -0.08 0.415 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.555 1.045 0.745 1.135 ;
        RECT 0.655 0.265 0.745 1.135 ;
        RECT 0.555 0.265 0.745 0.355 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.865 0.16 1.075 ;
      RECT 0.07 0.865 0.565 0.955 ;
      RECT 0.475 0.445 0.565 0.955 ;
      RECT 0.07 0.445 0.565 0.535 ;
      RECT 0.07 0.265 0.16 0.535 ;
  END
END BUFX3P5H7R

MACRO BUFX4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX4H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.835 0.855 0.925 1.48 ;
        RECT 0.325 1.07 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.835 -0.08 0.925 0.345 ;
        RECT 0.325 -0.08 0.415 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.165 0.625 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.555 1.045 0.745 1.135 ;
        RECT 0.655 0.265 0.745 1.135 ;
        RECT 0.555 0.265 0.745 0.355 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.075 0.865 0.165 1.035 ;
      RECT 0.075 0.865 0.549 0.955 ;
      RECT 0.459 0.445 0.549 0.955 ;
      RECT 0.075 0.445 0.549 0.535 ;
      RECT 0.075 0.305 0.165 0.535 ;
  END
END BUFX4H7R

MACRO BUFX5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX5H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.99 1.07 1.08 1.48 ;
        RECT 0.49 1.07 0.58 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.965 -0.08 1.105 0.305 ;
        RECT 0.465 -0.08 0.605 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.405 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.24 0.205 1.33 1.155 ;
        RECT 0.715 0.855 1.33 0.945 ;
        RECT 0.74 0.395 1.33 0.485 ;
        RECT 0.74 0.34 0.83 0.485 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.215 0.885 0.625 0.975 ;
      RECT 0.535 0.41 0.625 0.975 ;
      RECT 0.535 0.64 0.985 0.73 ;
      RECT 0.24 0.41 0.625 0.5 ;
      RECT 0.24 0.285 0.33 0.5 ;
  END
END BUFX5H7R

MACRO BUFX6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX6H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 0.82 1.07 0.91 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.545 -0.08 1.685 0.305 ;
        RECT 1.045 -0.08 1.185 0.305 ;
        RECT 0.57 -0.08 0.66 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.05 0.625 0.23 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.545 0.855 1.645 0.945 ;
        RECT 1.555 0.395 1.645 0.945 ;
        RECT 0.795 0.395 1.645 0.485 ;
        RECT 1.32 0.22 1.41 0.485 ;
        RECT 1.07 0.855 1.16 1.17 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.88 0.16 1.195 ;
      RECT 0.045 0.88 0.41 0.97 ;
      RECT 0.32 0.22 0.41 0.97 ;
      RECT 0.32 0.625 1.465 0.715 ;
  END
END BUFX6H7R

MACRO BUFX7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX7H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.57 1.055 1.66 1.48 ;
        RECT 1.07 1.07 1.16 1.48 ;
        RECT 0.57 1.07 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.57 -0.08 1.66 0.345 ;
        RECT 1.045 -0.08 1.185 0.305 ;
        RECT 0.57 -0.08 0.66 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.175 0.61 0.375 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.32 0.22 1.41 1.008 ;
        RECT 0.82 0.855 1.41 0.945 ;
        RECT 0.795 0.395 1.41 0.485 ;
        RECT 0.82 0.855 0.91 0.997 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.32 0.855 0.41 1.08 ;
      RECT 0.32 0.855 0.555 0.945 ;
      RECT 0.465 0.42 0.555 0.945 ;
      RECT 0.465 0.625 1.065 0.715 ;
      RECT 0.32 0.42 0.555 0.51 ;
      RECT 0.32 0.27 0.41 0.51 ;
  END
END BUFX7H7R

MACRO BUFX8H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX8H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.57 1.055 1.66 1.48 ;
        RECT 1.07 1.07 1.16 1.48 ;
        RECT 0.57 1.07 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.545 -0.08 1.685 0.305 ;
        RECT 1.045 -0.08 1.185 0.305 ;
        RECT 0.57 -0.08 0.66 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.05 0.625 0.23 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.82 0.855 1.91 0.945 ;
        RECT 1.82 0.205 1.91 0.945 ;
        RECT 0.795 0.395 1.91 0.485 ;
        RECT 1.32 0.855 1.41 1.17 ;
        RECT 1.32 0.22 1.41 0.485 ;
        RECT 0.82 0.855 0.91 1.195 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.32 0.205 0.41 1.09 ;
      RECT 0.32 0.625 1.665 0.715 ;
  END
END BUFX8H7R

MACRO DFFNQX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNQX1H7R 0 0 ;
  SIZE 4.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.6 1.48 ;
        RECT 4.319 1.022 4.459 1.48 ;
        RECT 3.474 1.24 3.614 1.48 ;
        RECT 2.227 1.156 2.367 1.48 ;
        RECT 1.37 1.225 1.51 1.48 ;
        RECT 0.31 1.15 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.6 0.08 ;
        RECT 4.294 -0.08 4.384 0.45 ;
        RECT 3.435 -0.08 3.525 0.41 ;
        RECT 2.227 -0.08 2.367 0.175 ;
        RECT 1.385 -0.08 1.525 0.16 ;
        RECT 0.325 -0.08 0.465 0.16 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.625 0.37 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.485 0.455 0.575 0.695 ;
        RECT 0.425 0.455 0.575 0.545 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.805 0.955 3.945 1.045 ;
        RECT 3.855 0.32 3.945 1.045 ;
        RECT 3.66 0.32 3.945 0.41 ;
      LAYER MET2 ;
        RECT 3.85 0.23 3.95 0.76 ;
      LAYER VIA1 ;
        RECT 3.855 0.455 3.945 0.545 ;
    END
  END Q
  OBS
    LAYER MET1 ;
      RECT 3.732 1.14 4.184 1.23 ;
      RECT 4.094 0.31 4.184 1.23 ;
      RECT 3.215 1.14 3.356 1.23 ;
      RECT 3.69 1.14 4.184 1.209 ;
      RECT 3.215 1.14 3.398 1.209 ;
      RECT 3.652 1.14 4.184 1.169 ;
      RECT 3.215 1.14 3.436 1.169 ;
      RECT 3.398 1.06 3.69 1.15 ;
      RECT 3.318 1.121 3.77 1.15 ;
      RECT 3.356 1.081 3.732 1.15 ;
      RECT 4.044 0.31 4.184 0.45 ;
      RECT 2.815 0.96 3.202 1.05 ;
      RECT 3.225 0.525 3.271 1.004 ;
      RECT 3.164 0.941 3.271 1.004 ;
      RECT 3.202 0.91 3.225 1.039 ;
      RECT 3.225 0.57 3.315 0.959 ;
      RECT 3.225 0.66 3.73 0.75 ;
      RECT 3.223 0.501 3.225 0.629 ;
      RECT 3.177 0.477 3.223 0.605 ;
      RECT 3.131 0.431 3.177 0.559 ;
      RECT 3.085 0.385 3.131 0.513 ;
      RECT 3.047 0.431 3.177 0.471 ;
      RECT 2.935 0.362 3.085 0.452 ;
      RECT 0.54 1.14 0.855 1.23 ;
      RECT 0.54 0.96 0.63 1.23 ;
      RECT 0.07 0.96 0.63 1.05 ;
      RECT 0.07 0.25 0.16 1.05 ;
      RECT 2.839 0.755 3.135 0.845 ;
      RECT 2.839 0.557 2.929 0.845 ;
      RECT 2.798 0.514 2.888 0.596 ;
      RECT 2.752 0.17 2.842 0.552 ;
      RECT 2.148 0.265 2.541 0.355 ;
      RECT 2.137 0.221 2.148 0.35 ;
      RECT 1.229 0.25 1.602 0.34 ;
      RECT 0.07 0.25 0.681 0.34 ;
      RECT 2.137 0.265 2.587 0.332 ;
      RECT 2.091 0.193 2.137 0.321 ;
      RECT 1.187 0.25 1.644 0.319 ;
      RECT 1.149 0.25 1.682 0.279 ;
      RECT 2.503 0.246 2.636 0.279 ;
      RECT 2.587 0.175 2.598 0.304 ;
      RECT 2.053 0.246 2.186 0.279 ;
      RECT 2.598 0.17 2.842 0.26 ;
      RECT 1.644 0.17 2.091 0.26 ;
      RECT 1.602 0.191 1.644 0.319 ;
      RECT 0.591 0.231 1.267 0.26 ;
      RECT 2.541 0.204 2.842 0.26 ;
      RECT 1.564 0.231 2.148 0.26 ;
      RECT 0.591 0.191 1.229 0.26 ;
      RECT 0.591 0.17 1.187 0.26 ;
      RECT 1.643 1.14 2.077 1.23 ;
      RECT 1.987 0.845 2.077 1.23 ;
      RECT 1.632 1.096 1.643 1.225 ;
      RECT 1.586 1.068 1.632 1.196 ;
      RECT 1.548 1.121 1.681 1.154 ;
      RECT 1.05 1.045 1.586 1.135 ;
      RECT 1.05 0.745 1.14 1.135 ;
      RECT 1.987 0.845 2.662 0.949 ;
      RECT 2.572 0.445 2.662 0.949 ;
      RECT 2.572 0.72 2.747 0.86 ;
      RECT 0.94 0.745 1.14 0.835 ;
      RECT 1.945 0.445 2.662 0.535 ;
      RECT 1.715 0.37 1.81 1.045 ;
      RECT 1.255 0.865 1.81 0.955 ;
      RECT 1.7 0.37 1.81 0.955 ;
      RECT 1.255 0.72 1.345 0.955 ;
      RECT 1.7 0.665 2.432 0.755 ;
      RECT 1.7 0.37 1.84 0.46 ;
      RECT 0.76 0.941 0.96 1.031 ;
      RECT 0.76 0.373 0.85 1.031 ;
      RECT 1.515 0.43 1.605 0.655 ;
      RECT 0.76 0.43 1.605 0.52 ;
      RECT 0.806 0.35 0.955 0.52 ;
  END
END DFFNQX1H7R

MACRO DFFNQX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNQX2H7R 0 0 ;
  SIZE 4.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.6 1.48 ;
        RECT 4.319 1.022 4.459 1.48 ;
        RECT 3.434 1.24 3.574 1.48 ;
        RECT 2.212 1.03 2.352 1.48 ;
        RECT 1.35 1.205 1.49 1.48 ;
        RECT 0.31 1.15 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.6 0.08 ;
        RECT 4.294 -0.08 4.384 0.45 ;
        RECT 3.395 -0.08 3.485 0.345 ;
        RECT 2.227 -0.08 2.367 0.175 ;
        RECT 1.376 -0.08 1.516 0.175 ;
        RECT 0.325 -0.08 0.465 0.16 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.625 0.37 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.485 0.455 0.575 0.695 ;
        RECT 0.425 0.455 0.575 0.545 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.855 0.38 3.945 0.965 ;
        RECT 3.62 0.38 3.945 0.47 ;
      LAYER MET2 ;
        RECT 3.85 0.23 3.95 0.76 ;
      LAYER VIA1 ;
        RECT 3.855 0.455 3.945 0.545 ;
    END
  END Q
  OBS
    LAYER MET1 ;
      RECT 3.175 1.14 3.315 1.23 ;
      RECT 3.175 1.14 3.357 1.209 ;
      RECT 3.175 1.14 3.395 1.169 ;
      RECT 4.094 0.31 4.184 1.15 ;
      RECT 3.277 1.121 4.184 1.15 ;
      RECT 3.357 1.06 4.184 1.15 ;
      RECT 3.315 1.081 4.184 1.15 ;
      RECT 4.044 0.31 4.184 0.45 ;
      RECT 2.815 0.96 3.207 1.05 ;
      RECT 3.225 0.43 3.271 1.009 ;
      RECT 3.225 0.475 3.315 0.964 ;
      RECT 3.169 0.941 3.315 0.964 ;
      RECT 3.207 0.913 3.225 1.041 ;
      RECT 3.225 0.612 3.69 0.702 ;
      RECT 3.18 0.384 3.225 0.513 ;
      RECT 3.142 0.43 3.271 0.471 ;
      RECT 2.885 0.362 3.18 0.452 ;
      RECT 0.54 1.14 0.828 1.23 ;
      RECT 0.54 0.96 0.63 1.23 ;
      RECT 0.07 0.96 0.63 1.05 ;
      RECT 0.07 0.25 0.16 1.05 ;
      RECT 3.031 0.755 3.135 0.845 ;
      RECT 1.292 0.275 1.544 0.365 ;
      RECT 2.186 0.265 2.438 0.355 ;
      RECT 0.07 0.25 0.681 0.34 ;
      RECT 2.571 0.17 2.705 0.26 ;
      RECT 1.687 0.17 2.053 0.26 ;
      RECT 0.591 0.17 1.149 0.26 ;
      RECT 2.993 0.736 3.031 0.845 ;
      RECT 2.979 0.71 2.993 0.838 ;
      RECT 2.933 0.68 2.979 0.808 ;
      RECT 2.887 0.634 2.933 0.762 ;
      RECT 2.841 0.588 2.887 0.716 ;
      RECT 2.795 0.542 2.841 0.67 ;
      RECT 2.751 0.17 2.795 0.625 ;
      RECT 2.705 0.17 2.751 0.58 ;
      RECT 2.533 0.17 2.571 0.279 ;
      RECT 2.522 0.175 2.533 0.304 ;
      RECT 2.476 0.204 2.522 0.332 ;
      RECT 2.438 0.246 2.476 0.355 ;
      RECT 2.148 0.246 2.186 0.355 ;
      RECT 2.137 0.221 2.148 0.35 ;
      RECT 2.091 0.193 2.137 0.321 ;
      RECT 2.053 0.17 2.091 0.279 ;
      RECT 1.649 0.17 1.687 0.279 ;
      RECT 1.628 0.18 1.649 0.309 ;
      RECT 1.582 0.214 1.628 0.342 ;
      RECT 1.544 0.256 1.582 0.365 ;
      RECT 1.254 0.256 1.292 0.365 ;
      RECT 1.233 0.226 1.254 0.355 ;
      RECT 1.187 0.193 1.233 0.321 ;
      RECT 1.149 0.17 1.187 0.279 ;
      RECT 1.643 1.14 2.077 1.23 ;
      RECT 1.987 0.845 2.077 1.23 ;
      RECT 1.612 1.086 1.643 1.215 ;
      RECT 1.566 1.048 1.612 1.176 ;
      RECT 1.566 1.121 1.681 1.176 ;
      RECT 1.528 1.025 1.566 1.134 ;
      RECT 1.02 1.025 1.566 1.115 ;
      RECT 1.02 0.745 1.11 1.115 ;
      RECT 1.987 0.845 2.615 0.935 ;
      RECT 2.525 0.445 2.615 0.935 ;
      RECT 2.525 0.745 2.75 0.835 ;
      RECT 0.91 0.745 1.11 0.835 ;
      RECT 1.945 0.445 2.615 0.535 ;
      RECT 1.715 0.364 1.805 1.045 ;
      RECT 1.256 0.76 1.805 0.85 ;
      RECT 1.256 0.695 1.346 0.85 ;
      RECT 1.715 0.665 2.432 0.755 ;
      RECT 0.73 0.941 0.93 1.031 ;
      RECT 0.73 0.398 0.82 1.031 ;
      RECT 1.516 0.455 1.606 0.67 ;
      RECT 0.73 0.455 1.606 0.545 ;
      RECT 0.801 0.35 0.955 0.545 ;
      RECT 0.776 0.362 0.955 0.545 ;
  END
END DFFNQX2H7R

MACRO DFFNQX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNQX3H7R 0 0 ;
  SIZE 4.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.8 1.48 ;
        RECT 4.614 0.905 4.704 1.48 ;
        RECT 4.094 1.215 4.234 1.48 ;
        RECT 3.484 1.24 3.624 1.48 ;
        RECT 2.202 1.156 2.342 1.48 ;
        RECT 1.37 1.225 1.51 1.48 ;
        RECT 0.31 1.15 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.8 0.08 ;
        RECT 4.564 -0.08 4.654 0.45 ;
        RECT 3.951 -0.08 4.091 0.205 ;
        RECT 3.421 -0.08 3.561 0.37 ;
        RECT 2.202 -0.08 2.342 0.175 ;
        RECT 1.38 -0.08 1.52 0.175 ;
        RECT 0.325 -0.08 0.465 0.16 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.625 0.37 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.485 0.455 0.575 0.695 ;
        RECT 0.425 0.455 0.575 0.545 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.814 0.855 4.175 0.945 ;
        RECT 4.076 0.32 4.175 0.945 ;
        RECT 3.686 0.32 4.175 0.41 ;
      LAYER MET2 ;
        RECT 4.05 0.63 4.15 1.16 ;
      LAYER VIA1 ;
        RECT 4.055 0.855 4.145 0.945 ;
    END
  END Q
  OBS
    LAYER MET1 ;
      RECT 3.226 1.14 3.366 1.23 ;
      RECT 3.226 1.14 3.412 1.207 ;
      RECT 3.328 1.121 3.471 1.144 ;
      RECT 3.412 1.045 3.433 1.174 ;
      RECT 4.364 0.31 4.454 1.125 ;
      RECT 3.366 1.079 4.454 1.125 ;
      RECT 3.433 1.035 4.454 1.125 ;
      RECT 4.314 0.31 4.454 0.45 ;
      RECT 2.79 0.96 3.242 1.05 ;
      RECT 3.281 0.511 3.327 0.988 ;
      RECT 3.204 0.941 3.327 0.988 ;
      RECT 3.242 0.902 3.281 1.031 ;
      RECT 3.281 0.556 3.371 0.943 ;
      RECT 3.281 0.612 3.956 0.702 ;
      RECT 3.247 0.471 3.281 0.599 ;
      RECT 3.201 0.431 3.247 0.559 ;
      RECT 3.155 0.385 3.201 0.513 ;
      RECT 3.117 0.362 3.155 0.471 ;
      RECT 2.946 0.362 3.155 0.452 ;
      RECT 0.54 1.14 0.828 1.23 ;
      RECT 0.54 0.96 0.63 1.23 ;
      RECT 0.07 0.96 0.63 1.05 ;
      RECT 0.07 0.25 0.16 1.05 ;
      RECT 2.904 0.755 3.11 0.845 ;
      RECT 2.814 0.17 2.817 0.845 ;
      RECT 1.292 0.275 1.548 0.365 ;
      RECT 2.161 0.265 2.478 0.355 ;
      RECT 0.07 0.25 0.681 0.34 ;
      RECT 2.611 0.17 2.727 0.26 ;
      RECT 1.691 0.17 2.028 0.26 ;
      RECT 0.591 0.17 1.149 0.26 ;
      RECT 2.863 0.557 2.904 0.845 ;
      RECT 2.817 0.514 2.863 0.845 ;
      RECT 2.773 0.17 2.814 0.596 ;
      RECT 2.727 0.17 2.773 0.552 ;
      RECT 2.573 0.17 2.611 0.279 ;
      RECT 2.562 0.175 2.573 0.304 ;
      RECT 2.516 0.204 2.562 0.332 ;
      RECT 2.478 0.246 2.516 0.355 ;
      RECT 2.123 0.246 2.161 0.355 ;
      RECT 2.082 0.206 2.123 0.335 ;
      RECT 2.074 0.17 2.082 0.31 ;
      RECT 2.028 0.17 2.074 0.283 ;
      RECT 1.653 0.17 1.691 0.279 ;
      RECT 1.632 0.18 1.653 0.309 ;
      RECT 1.586 0.214 1.632 0.342 ;
      RECT 1.548 0.256 1.586 0.365 ;
      RECT 1.254 0.256 1.292 0.365 ;
      RECT 1.233 0.226 1.254 0.355 ;
      RECT 1.187 0.193 1.233 0.321 ;
      RECT 1.149 0.17 1.187 0.279 ;
      RECT 1.643 1.14 2.052 1.23 ;
      RECT 1.962 0.845 2.052 1.23 ;
      RECT 1.632 1.096 1.643 1.225 ;
      RECT 1.586 1.068 1.632 1.196 ;
      RECT 1.548 1.121 1.681 1.154 ;
      RECT 1.02 1.045 1.586 1.135 ;
      RECT 1.02 0.745 1.11 1.135 ;
      RECT 1.962 0.845 2.637 0.949 ;
      RECT 2.547 0.445 2.637 0.949 ;
      RECT 2.547 0.72 2.699 0.86 ;
      RECT 0.91 0.745 1.11 0.835 ;
      RECT 1.92 0.445 2.637 0.535 ;
      RECT 1.715 0.364 1.805 1.045 ;
      RECT 1.256 0.755 1.805 0.845 ;
      RECT 1.715 0.665 2.432 0.755 ;
      RECT 1.256 0.695 1.346 0.845 ;
      RECT 0.73 0.941 0.93 1.031 ;
      RECT 0.73 0.398 0.82 1.031 ;
      RECT 1.516 0.455 1.606 0.665 ;
      RECT 0.73 0.455 1.606 0.545 ;
      RECT 0.801 0.35 0.955 0.545 ;
      RECT 0.776 0.362 0.955 0.545 ;
  END
END DFFNQX3H7R

MACRO DFFNRX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNRX0P5H7R 0 0 ;
  SIZE 6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6 1.48 ;
        RECT 5.53 1.225 5.67 1.48 ;
        RECT 5.02 1.225 5.16 1.48 ;
        RECT 3.734 1.188 3.874 1.48 ;
        RECT 1.756 1.225 1.896 1.48 ;
        RECT 0.815 1.14 0.905 1.48 ;
        RECT 0.32 1.035 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6 0.08 ;
        RECT 5.558 -0.08 5.648 0.375 ;
        RECT 5.03 -0.08 5.12 0.36 ;
        RECT 3.675 -0.08 3.815 0.175 ;
        RECT 2.252 -0.08 2.342 0.44 ;
        RECT 1.642 -0.08 1.782 0.235 ;
        RECT 0.815 -0.08 0.905 0.35 ;
        RECT 0.32 -0.08 0.41 0.365 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 5.655 0.49 5.745 0.79 ;
      LAYER MET2 ;
        RECT 5.65 0.425 5.75 0.96 ;
      LAYER VIA1 ;
        RECT 5.655 0.655 5.745 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.905 0.655 5.175 0.755 ;
      LAYER MET2 ;
        RECT 5.05 0.43 5.15 0.96 ;
      LAYER VIA1 ;
        RECT 5.055 0.655 5.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.905 0.175 1.045 ;
        RECT 0.055 0.275 0.175 0.415 ;
        RECT 0.055 0.275 0.145 1.045 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.78 1.21 0.87 ;
        RECT 1.055 0.257 1.2 0.347 ;
        RECT 1.055 0.257 1.145 0.87 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.481 1.467 0.585 ;
        RECT 1.255 0.425 1.345 0.585 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END RN
  OBS
    LAYER MET1 ;
      RECT 4.048 1.12 4.785 1.21 ;
      RECT 4.695 0.745 4.785 1.21 ;
      RECT 4.018 1.067 4.048 1.195 ;
      RECT 3.972 1.029 4.018 1.157 ;
      RECT 5.475 0.72 5.565 1.135 ;
      RECT 4.695 1.045 5.565 1.135 ;
      RECT 3.972 1.101 4.086 1.157 ;
      RECT 3.926 0.983 3.972 1.111 ;
      RECT 3.888 0.96 3.926 1.069 ;
      RECT 2.741 0.96 3.926 1.05 ;
      RECT 5.84 0.299 5.93 1.045 ;
      RECT 5.475 0.955 5.93 1.045 ;
      RECT 3.157 0.589 3.247 1.05 ;
      RECT 2.741 0.766 2.831 1.05 ;
      RECT 2.511 0.766 2.831 0.856 ;
      RECT 4.211 0.745 4.785 0.835 ;
      RECT 2.511 0.716 2.601 0.856 ;
      RECT 4.211 0.546 4.301 0.835 ;
      RECT 4.161 0.546 4.301 0.636 ;
      RECT 5.275 0.299 5.365 0.955 ;
      RECT 4.585 0.17 4.675 0.63 ;
      RECT 2.617 0.51 2.761 0.6 ;
      RECT 2.617 0.51 2.807 0.577 ;
      RECT 4.585 0.45 5.365 0.54 ;
      RECT 2.723 0.491 2.853 0.531 ;
      RECT 2.761 0.449 2.853 0.531 ;
      RECT 2.807 0.403 2.899 0.485 ;
      RECT 2.853 0.357 2.945 0.439 ;
      RECT 2.899 0.311 2.991 0.393 ;
      RECT 3.599 0.265 3.914 0.355 ;
      RECT 3.588 0.221 3.599 0.35 ;
      RECT 3.588 0.265 3.96 0.332 ;
      RECT 3.542 0.193 3.588 0.321 ;
      RECT 3.037 0.183 3.063 0.311 ;
      RECT 2.945 0.265 3.063 0.311 ;
      RECT 2.991 0.219 3.037 0.347 ;
      RECT 3.063 0.17 3.101 0.279 ;
      RECT 3.876 0.246 4.009 0.279 ;
      RECT 3.96 0.175 3.971 0.304 ;
      RECT 3.504 0.246 3.637 0.279 ;
      RECT 3.971 0.17 4.675 0.26 ;
      RECT 3.063 0.17 3.542 0.26 ;
      RECT 3.914 0.204 4.675 0.26 ;
      RECT 4.145 0.94 4.574 1.03 ;
      RECT 4.135 0.897 4.145 1.025 ;
      RECT 4.089 0.869 4.135 0.997 ;
      RECT 4.043 0.823 4.089 0.951 ;
      RECT 4.043 0.921 4.183 0.951 ;
      RECT 3.999 0.418 4.043 0.906 ;
      RECT 3.953 0.463 4.043 0.861 ;
      RECT 3.95 0.823 4.089 0.837 ;
      RECT 3.395 0.745 4.043 0.835 ;
      RECT 4.089 0.35 4.135 0.463 ;
      RECT 4.043 0.373 4.089 0.509 ;
      RECT 4.089 0.35 4.49 0.44 ;
      RECT 2.921 0.78 3.061 0.87 ;
      RECT 2.921 0.546 3.011 0.87 ;
      RECT 3.355 0.52 3.78 0.61 ;
      RECT 2.967 0.501 3.057 0.584 ;
      RECT 3.355 0.35 3.445 0.61 ;
      RECT 3.011 0.456 3.103 0.538 ;
      RECT 3.057 0.41 3.178 0.459 ;
      RECT 3.103 0.368 3.14 0.497 ;
      RECT 3.14 0.35 3.445 0.44 ;
      RECT 1.003 1.14 1.623 1.23 ;
      RECT 1.003 1.14 1.669 1.207 ;
      RECT 1.585 1.121 1.715 1.161 ;
      RECT 1.623 1.079 1.715 1.161 ;
      RECT 1.623 1.079 1.761 1.115 ;
      RECT 1.669 1.033 1.779 1.083 ;
      RECT 1.669 1.033 1.817 1.055 ;
      RECT 1.779 0.946 2.651 1.036 ;
      RECT 1.715 0.987 2.651 1.036 ;
      RECT 1.761 0.955 1.779 1.083 ;
      RECT 2.331 0.53 2.421 1.036 ;
      RECT 2.168 0.53 2.527 0.62 ;
      RECT 2.437 0.17 2.527 0.62 ;
      RECT 2.134 0.475 2.168 0.603 ;
      RECT 2.088 0.435 2.134 0.563 ;
      RECT 2.088 0.511 2.206 0.563 ;
      RECT 2.042 0.389 2.088 0.517 ;
      RECT 1.998 0.255 2.042 0.472 ;
      RECT 1.952 0.255 2.042 0.427 ;
      RECT 2.437 0.17 2.842 0.26 ;
      RECT 0.55 0.96 1.518 1.05 ;
      RECT 0.55 0.96 1.564 1.027 ;
      RECT 1.48 0.941 1.61 0.981 ;
      RECT 0.55 0.27 0.64 1.05 ;
      RECT 1.518 0.899 1.61 0.981 ;
      RECT 1.564 0.853 1.656 0.935 ;
      RECT 1.564 0.853 1.702 0.889 ;
      RECT 1.61 0.807 1.72 0.857 ;
      RECT 1.61 0.807 1.758 0.829 ;
      RECT 1.72 0.72 2.241 0.81 ;
      RECT 1.656 0.761 2.241 0.81 ;
      RECT 1.702 0.729 1.72 0.857 ;
      RECT 0.235 0.625 0.64 0.715 ;
      RECT 1.302 0.78 1.442 0.87 ;
      RECT 1.302 0.78 1.488 0.847 ;
      RECT 1.404 0.761 1.534 0.801 ;
      RECT 1.442 0.719 1.557 0.767 ;
      RECT 1.557 0.304 1.603 0.732 ;
      RECT 1.488 0.673 1.603 0.732 ;
      RECT 1.534 0.638 1.557 0.767 ;
      RECT 1.557 0.349 1.647 0.687 ;
      RECT 1.557 0.53 1.907 0.62 ;
      RECT 1.526 0.265 1.557 0.394 ;
      RECT 1.488 0.25 1.526 0.359 ;
      RECT 1.377 0.25 1.526 0.34 ;
      RECT 2.036 1.14 3.617 1.23 ;
  END
END DFFNRX0P5H7R

MACRO DFFNRX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNRX1H7R 0 0 ;
  SIZE 7 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7 1.48 ;
        RECT 6.495 1.195 6.635 1.48 ;
        RECT 5.71 1.225 5.85 1.48 ;
        RECT 4.43 1.225 4.57 1.48 ;
        RECT 2.225 0.89 2.315 1.48 ;
        RECT 0.805 1.195 0.945 1.48 ;
        RECT 0.335 1.195 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7 0.08 ;
        RECT 6.505 -0.08 6.595 0.345 ;
        RECT 6.015 -0.08 6.105 0.365 ;
        RECT 5.21 -0.08 5.3 0.365 ;
        RECT 4.43 -0.08 4.57 0.175 ;
        RECT 1.975 -0.08 2.065 0.38 ;
        RECT 0.845 -0.08 0.935 0.36 ;
        RECT 0.32 -0.08 0.41 0.335 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.35 0.695 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.82 0.625 1.045 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.792 0.425 6.945 0.575 ;
        RECT 6.792 0.31 6.882 0.925 ;
      LAYER MET2 ;
        RECT 6.85 0.23 6.95 0.76 ;
      LAYER VIA1 ;
        RECT 6.855 0.455 6.945 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.255 0.31 6.345 0.925 ;
      LAYER MET2 ;
        RECT 6.25 0.425 6.35 0.96 ;
      LAYER VIA1 ;
        RECT 6.255 0.655 6.345 0.745 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.705 0.455 3.795 0.87 ;
        RECT 3.625 0.455 3.795 0.545 ;
      LAYER MET2 ;
        RECT 3.65 0.23 3.75 0.76 ;
      LAYER VIA1 ;
        RECT 3.655 0.455 3.745 0.545 ;
    END
  END RN
  OBS
    LAYER MET1 ;
      RECT 6.015 1.015 6.68 1.105 ;
      RECT 6.59 0.575 6.68 1.105 ;
      RECT 6.015 0.561 6.105 1.105 ;
      RECT 5.972 0.471 6.015 0.6 ;
      RECT 5.972 0.516 6.061 0.6 ;
      RECT 5.926 0.427 5.972 0.555 ;
      RECT 5.88 0.381 5.926 0.509 ;
      RECT 5.835 0.305 5.88 0.464 ;
      RECT 5.789 0.381 5.926 0.418 ;
      RECT 5.415 0.305 5.88 0.395 ;
      RECT 5.05 1.045 5.14 1.23 ;
      RECT 5.05 1.045 5.905 1.135 ;
      RECT 5.815 0.629 5.905 1.135 ;
      RECT 3.445 0.78 3.59 0.87 ;
      RECT 3.445 0.17 3.535 0.87 ;
      RECT 5.785 0.546 5.815 0.674 ;
      RECT 5.739 0.508 5.785 0.636 ;
      RECT 5.739 0.584 5.861 0.636 ;
      RECT 5.701 0.485 5.739 0.594 ;
      RECT 4.951 0.485 5.739 0.575 ;
      RECT 4.951 0.265 5.041 0.575 ;
      RECT 4.354 0.265 5.041 0.355 ;
      RECT 4.343 0.221 4.354 0.35 ;
      RECT 4.297 0.193 4.343 0.321 ;
      RECT 4.259 0.246 4.392 0.279 ;
      RECT 3.445 0.17 4.297 0.26 ;
      RECT 2.855 0.96 4.156 1.05 ;
      RECT 2.855 0.96 4.202 1.027 ;
      RECT 4.118 0.941 4.251 0.974 ;
      RECT 4.202 0.87 4.213 0.999 ;
      RECT 2.855 0.93 2.995 1.05 ;
      RECT 5.5 0.835 5.64 0.955 ;
      RECT 4.156 0.899 5.64 0.955 ;
      RECT 4.213 0.865 5.64 0.955 ;
      RECT 4.242 0.665 5.25 0.755 ;
      RECT 4.22 0.616 4.242 0.744 ;
      RECT 4.182 0.665 5.25 0.714 ;
      RECT 4.08 0.605 4.22 0.695 ;
      RECT 4.08 0.646 4.28 0.695 ;
      RECT 2.44 1.14 4.236 1.23 ;
      RECT 2.44 1.14 4.282 1.207 ;
      RECT 4.85 1.045 4.94 1.195 ;
      RECT 4.198 1.121 4.331 1.154 ;
      RECT 4.282 1.05 4.293 1.179 ;
      RECT 4.293 1.045 4.94 1.135 ;
      RECT 4.236 1.079 4.94 1.135 ;
      RECT 3.9 0.78 4.05 0.87 ;
      RECT 3.9 0.486 3.99 0.87 ;
      RECT 4.524 0.445 4.665 0.575 ;
      RECT 4.277 0.445 4.665 0.535 ;
      RECT 3.9 0.486 4.036 0.524 ;
      RECT 4.231 0.383 4.277 0.511 ;
      RECT 3.946 0.441 4.049 0.495 ;
      RECT 4.193 0.445 4.665 0.469 ;
      RECT 3.946 0.441 4.087 0.469 ;
      RECT 4.049 0.36 4.231 0.45 ;
      RECT 4.277 0.426 4.316 0.535 ;
      RECT 4.036 0.366 4.049 0.495 ;
      RECT 3.99 0.406 4.278 0.45 ;
      RECT 3.99 0.396 4.277 0.45 ;
      RECT 3.14 0.78 3.285 0.87 ;
      RECT 3.195 0.275 3.285 0.87 ;
      RECT 2.405 0.495 3.285 0.585 ;
      RECT 2.405 0.29 2.495 0.585 ;
      RECT 2.2 0.29 2.495 0.38 ;
      RECT 1.035 1.14 2.135 1.23 ;
      RECT 2.045 0.7 2.135 1.23 ;
      RECT 0.515 1.015 0.655 1.21 ;
      RECT 1.035 1.015 1.125 1.23 ;
      RECT 0.07 1.015 1.125 1.105 ;
      RECT 0.07 0.26 0.16 1.105 ;
      RECT 2.96 0.675 3.05 0.815 ;
      RECT 2.045 0.7 3.05 0.79 ;
      RECT 2.63 0.88 2.72 1.045 ;
      RECT 2.405 0.88 2.72 0.97 ;
      RECT 1.435 0.935 1.955 1.025 ;
      RECT 1.865 0.52 1.955 1.025 ;
      RECT 1.435 0.35 1.525 1.025 ;
      RECT 1.865 0.52 2.27 0.61 ;
      RECT 1.385 0.35 1.525 0.44 ;
      RECT 0.6 0.835 1.295 0.925 ;
      RECT 1.205 0.17 1.295 0.925 ;
      RECT 1.685 0.17 1.775 0.845 ;
      RECT 0.6 0.26 0.69 0.925 ;
      RECT 1.205 0.17 1.775 0.26 ;
  END
END DFFNRX1H7R

MACRO DFFNRX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNRX2H7R 0 0 ;
  SIZE 7 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7 1.48 ;
        RECT 6.439 1.07 6.529 1.48 ;
        RECT 5.61 1.225 5.75 1.48 ;
        RECT 4.36 1.225 4.5 1.48 ;
        RECT 2.215 0.89 2.305 1.48 ;
        RECT 0.81 1.225 0.95 1.48 ;
        RECT 0.335 1.11 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7 0.08 ;
        RECT 6.825 -0.08 6.915 0.33 ;
        RECT 6.325 -0.08 6.415 0.33 ;
        RECT 5.845 -0.08 5.935 0.36 ;
        RECT 5.125 -0.08 5.215 0.365 ;
        RECT 4.36 -0.08 4.505 0.175 ;
        RECT 1.965 -0.08 2.055 0.36 ;
        RECT 0.84 -0.08 0.93 0.36 ;
        RECT 0.32 -0.08 0.41 0.335 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.35 0.695 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.625 1.035 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.655 0.83 6.805 0.92 ;
        RECT 6.655 0.425 6.745 0.92 ;
        RECT 6.575 0.21 6.665 0.515 ;
      LAYER MET2 ;
        RECT 6.65 0.425 6.75 0.96 ;
      LAYER VIA1 ;
        RECT 6.655 0.655 6.745 0.745 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.105 0.455 6.195 0.93 ;
        RECT 6.075 0.335 6.165 0.545 ;
        RECT 6.025 0.455 6.195 0.545 ;
      LAYER MET2 ;
        RECT 6.05 0.23 6.15 0.76 ;
      LAYER VIA1 ;
        RECT 6.055 0.455 6.145 0.545 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.655 0.35 3.805 0.44 ;
        RECT 3.655 0.35 3.745 0.59 ;
      LAYER MET2 ;
        RECT 3.65 0.23 3.75 0.76 ;
      LAYER VIA1 ;
        RECT 3.655 0.455 3.745 0.545 ;
    END
  END RN
  OBS
    LAYER MET1 ;
      RECT 5.845 1.06 6.231 1.15 ;
      RECT 5.845 1.06 6.277 1.127 ;
      RECT 6.193 1.041 6.323 1.081 ;
      RECT 5.845 0.558 5.935 1.15 ;
      RECT 6.231 0.999 6.323 1.081 ;
      RECT 6.277 0.953 6.369 1.035 ;
      RECT 6.323 0.907 6.415 0.989 ;
      RECT 6.323 0.907 6.461 0.943 ;
      RECT 6.369 0.861 6.465 0.918 ;
      RECT 6.415 0.815 6.511 0.893 ;
      RECT 6.461 0.79 6.465 0.918 ;
      RECT 6.465 0.62 6.555 0.848 ;
      RECT 5.844 0.489 5.845 0.618 ;
      RECT 5.798 0.466 5.844 0.594 ;
      RECT 5.798 0.513 5.891 0.594 ;
      RECT 5.752 0.42 5.798 0.548 ;
      RECT 5.706 0.374 5.752 0.502 ;
      RECT 5.66 0.328 5.706 0.456 ;
      RECT 5.622 0.374 5.752 0.414 ;
      RECT 5.32 0.305 5.66 0.395 ;
      RECT 4.98 1.045 5.07 1.185 ;
      RECT 4.98 1.045 5.755 1.135 ;
      RECT 5.665 0.634 5.755 1.135 ;
      RECT 3.44 0.78 3.585 0.87 ;
      RECT 3.44 0.17 3.53 0.87 ;
      RECT 5.63 0.548 5.665 0.677 ;
      RECT 5.584 0.508 5.63 0.636 ;
      RECT 5.584 0.589 5.711 0.636 ;
      RECT 5.546 0.485 5.584 0.594 ;
      RECT 4.904 0.485 5.584 0.575 ;
      RECT 4.904 0.265 4.994 0.575 ;
      RECT 4.284 0.265 4.994 0.355 ;
      RECT 4.273 0.221 4.284 0.35 ;
      RECT 4.227 0.193 4.273 0.321 ;
      RECT 4.189 0.246 4.322 0.279 ;
      RECT 3.44 0.17 4.227 0.26 ;
      RECT 2.845 0.96 4.059 1.05 ;
      RECT 2.845 0.96 4.105 1.027 ;
      RECT 4.021 0.941 4.154 0.967 ;
      RECT 4.105 0.863 4.131 0.991 ;
      RECT 4.131 0.85 5.57 0.955 ;
      RECT 4.059 0.899 5.57 0.955 ;
      RECT 4.04 0.665 5.18 0.755 ;
      RECT 4.04 0.595 4.13 0.755 ;
      RECT 2.395 1.14 4.149 1.23 ;
      RECT 2.395 1.14 4.195 1.207 ;
      RECT 4.78 1.045 4.87 1.195 ;
      RECT 4.111 1.121 4.244 1.154 ;
      RECT 4.195 1.05 4.206 1.179 ;
      RECT 4.206 1.045 4.87 1.135 ;
      RECT 4.149 1.079 4.87 1.135 ;
      RECT 3.71 0.78 3.925 0.87 ;
      RECT 3.835 0.519 3.925 0.87 ;
      RECT 4.248 0.485 4.605 0.575 ;
      RECT 4.202 0.424 4.248 0.552 ;
      RECT 3.881 0.474 3.971 0.557 ;
      RECT 4.156 0.378 4.202 0.506 ;
      RECT 4.156 0.466 4.286 0.506 ;
      RECT 3.925 0.429 4.015 0.512 ;
      RECT 3.925 0.429 4.06 0.468 ;
      RECT 4.118 0.424 4.248 0.464 ;
      RECT 4.015 0.355 4.156 0.445 ;
      RECT 3.971 0.384 4.015 0.512 ;
      RECT 3.13 0.78 3.28 0.87 ;
      RECT 3.19 0.29 3.28 0.87 ;
      RECT 2.42 0.29 2.51 0.61 ;
      RECT 2.19 0.29 3.28 0.38 ;
      RECT 1.2 1.14 2.125 1.23 ;
      RECT 2.035 0.7 2.125 1.23 ;
      RECT 1.2 1.045 1.29 1.23 ;
      RECT 0.581 1.045 1.29 1.135 ;
      RECT 0.57 1.001 0.581 1.13 ;
      RECT 0.526 1.045 1.29 1.102 ;
      RECT 0.48 0.57 0.57 1.057 ;
      RECT 0.48 1.026 0.619 1.057 ;
      RECT 0.451 1.001 0.581 1.02 ;
      RECT 0.07 0.915 0.57 1.005 ;
      RECT 0.07 0.3 0.16 1.005 ;
      RECT 2.035 0.7 3.04 0.79 ;
      RECT 2.95 0.65 3.04 0.79 ;
      RECT 1.38 0.935 1.945 1.025 ;
      RECT 1.855 0.52 1.945 1.025 ;
      RECT 1.38 0.35 1.47 1.025 ;
      RECT 1.855 0.52 2.26 0.61 ;
      RECT 1.38 0.35 1.52 0.44 ;
      RECT 0.66 0.865 1.29 0.955 ;
      RECT 1.2 0.17 1.29 0.955 ;
      RECT 0.66 0.325 0.75 0.955 ;
      RECT 1.675 0.17 1.765 0.845 ;
      RECT 0.575 0.325 0.75 0.415 ;
      RECT 1.2 0.17 1.765 0.26 ;
      RECT 2.395 0.88 2.735 0.98 ;
  END
END DFFNRX2H7R

MACRO DFFNRX4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNRX4H7R 0 0 ;
  SIZE 8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 8 1.48 ;
        RECT 7.393 1.025 7.533 1.48 ;
        RECT 6.833 0.845 6.923 1.48 ;
        RECT 6.183 1.225 6.323 1.48 ;
        RECT 5.673 1.225 5.813 1.48 ;
        RECT 4.415 1.225 4.555 1.48 ;
        RECT 2.23 0.89 2.32 1.48 ;
        RECT 0.81 1.225 0.95 1.48 ;
        RECT 0.335 1.2 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 8 0.08 ;
        RECT 7.433 -0.08 7.573 0.32 ;
        RECT 6.933 -0.08 7.073 0.32 ;
        RECT 6.433 -0.08 6.573 0.32 ;
        RECT 5.953 -0.08 6.093 0.34 ;
        RECT 5.285 -0.08 5.428 0.175 ;
        RECT 4.425 -0.08 4.57 0.175 ;
        RECT 1.895 0.285 2.21 0.375 ;
        RECT 1.895 -0.08 1.985 0.4 ;
        RECT 0.85 -0.08 0.94 0.345 ;
        RECT 0.32 -0.08 0.41 0.335 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.51 0.35 0.78 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.57 0.99 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.708 0.231 7.798 0.5 ;
        RECT 7.208 0.41 7.798 0.5 ;
        RECT 7.153 0.845 7.625 0.935 ;
        RECT 7.535 0.41 7.625 0.935 ;
        RECT 7.208 0.224 7.298 0.5 ;
        RECT 7.153 0.845 7.243 1.185 ;
        RECT 7.055 0.415 7.243 0.575 ;
      LAYER MET2 ;
        RECT 7.05 0.23 7.15 0.76 ;
      LAYER VIA1 ;
        RECT 7.055 0.455 7.145 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.208 0.41 6.798 0.5 ;
        RECT 6.708 0.23 6.798 0.5 ;
        RECT 6.455 0.41 6.563 0.905 ;
        RECT 6.208 0.235 6.298 0.5 ;
      LAYER MET2 ;
        RECT 6.45 0.425 6.55 0.96 ;
      LAYER VIA1 ;
        RECT 6.455 0.655 6.545 0.745 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.655 0.35 3.825 0.575 ;
      LAYER MET2 ;
        RECT 3.65 0.23 3.75 0.76 ;
      LAYER VIA1 ;
        RECT 3.655 0.455 3.745 0.545 ;
    END
  END RN
  OBS
    LAYER MET1 ;
      RECT 5.978 0.611 6.068 1.175 ;
      RECT 5.978 1.045 6.743 1.135 ;
      RECT 6.653 0.665 6.743 1.135 ;
      RECT 6.653 0.665 7.423 0.755 ;
      RECT 7.333 0.595 7.423 0.755 ;
      RECT 5.956 0.532 5.978 0.66 ;
      RECT 5.91 0.498 5.956 0.626 ;
      RECT 5.91 0.566 6.024 0.626 ;
      RECT 5.864 0.452 5.91 0.58 ;
      RECT 5.818 0.406 5.864 0.534 ;
      RECT 5.788 0.452 5.91 0.496 ;
      RECT 5.742 0.17 5.818 0.458 ;
      RECT 5.728 0.17 5.818 0.435 ;
      RECT 5.518 0.17 5.818 0.26 ;
      RECT 5.045 1.045 5.135 1.23 ;
      RECT 5.045 1.045 5.818 1.135 ;
      RECT 5.728 0.64 5.818 1.135 ;
      RECT 3.45 0.78 3.6 0.87 ;
      RECT 3.475 0.17 3.565 0.87 ;
      RECT 5.512 0.64 5.818 0.73 ;
      RECT 5.512 0.494 5.602 0.73 ;
      RECT 5.324 0.494 5.602 0.584 ;
      RECT 5.324 0.265 5.414 0.584 ;
      RECT 4.349 0.265 5.414 0.355 ;
      RECT 4.338 0.221 4.349 0.35 ;
      RECT 4.292 0.193 4.338 0.321 ;
      RECT 4.254 0.246 4.387 0.279 ;
      RECT 2.875 0.17 4.292 0.26 ;
      RECT 2.86 0.96 4.199 1.05 ;
      RECT 2.86 0.96 4.245 1.027 ;
      RECT 4.161 0.941 4.294 0.974 ;
      RECT 4.245 0.87 4.256 0.999 ;
      RECT 2.86 0.93 3 1.05 ;
      RECT 5.495 0.835 5.635 0.955 ;
      RECT 4.199 0.899 5.635 0.955 ;
      RECT 4.256 0.865 5.635 0.955 ;
      RECT 4.225 0.665 5.245 0.755 ;
      RECT 4.218 0.623 4.225 0.752 ;
      RECT 4.205 0.665 5.245 0.742 ;
      RECT 4.095 0.62 4.218 0.735 ;
      RECT 4.095 0.646 4.263 0.735 ;
      RECT 4.095 0.595 4.185 0.735 ;
      RECT 2.445 1.14 4.279 1.23 ;
      RECT 2.445 1.14 4.325 1.207 ;
      RECT 4.845 1.045 4.935 1.195 ;
      RECT 4.241 1.121 4.374 1.154 ;
      RECT 4.325 1.05 4.336 1.179 ;
      RECT 4.336 1.045 4.935 1.135 ;
      RECT 4.279 1.079 4.935 1.135 ;
      RECT 3.73 0.78 4.005 0.87 ;
      RECT 3.915 0.434 4.005 0.87 ;
      RECT 4.564 0.449 4.704 0.575 ;
      RECT 4.277 0.449 4.704 0.539 ;
      RECT 4.267 0.406 4.277 0.534 ;
      RECT 4.221 0.378 4.267 0.506 ;
      RECT 3.915 0.434 4.055 0.464 ;
      RECT 4.183 0.43 4.315 0.464 ;
      RECT 4.017 0.355 4.221 0.445 ;
      RECT 4.005 0.361 4.017 0.489 ;
      RECT 3.961 0.389 4.005 0.87 ;
      RECT 3.145 0.78 3.295 0.87 ;
      RECT 3.205 0.35 3.295 0.87 ;
      RECT 2.475 0.35 2.615 0.61 ;
      RECT 2.475 0.35 3.295 0.44 ;
      RECT 2.365 0.32 2.59 0.41 ;
      RECT 1.04 1.14 2.14 1.23 ;
      RECT 2.05 0.7 2.14 1.23 ;
      RECT 1.04 1.045 1.13 1.23 ;
      RECT 0.58 1.045 1.13 1.135 ;
      RECT 0.57 1.002 0.58 1.13 ;
      RECT 0.526 1.045 1.13 1.103 ;
      RECT 0.48 0.55 0.57 1.058 ;
      RECT 0.48 1.026 0.618 1.058 ;
      RECT 0.07 0.87 0.57 0.96 ;
      RECT 0.07 0.3 0.16 0.96 ;
      RECT 2.05 0.7 2.945 0.79 ;
      RECT 2.855 0.54 2.945 0.79 ;
      RECT 2.855 0.54 3.11 0.63 ;
      RECT 2.495 0.945 2.75 1.035 ;
      RECT 2.41 0.88 2.585 0.97 ;
      RECT 1.44 0.935 1.96 1.025 ;
      RECT 1.87 0.52 1.96 1.025 ;
      RECT 1.44 0.35 1.53 1.025 ;
      RECT 1.87 0.52 2.275 0.61 ;
      RECT 1.39 0.35 1.53 0.44 ;
      RECT 0.66 0.865 1.3 0.955 ;
      RECT 1.21 0.17 1.3 0.955 ;
      RECT 0.66 0.325 0.75 0.955 ;
      RECT 1.69 0.17 1.78 0.845 ;
      RECT 0.575 0.325 0.75 0.415 ;
      RECT 1.21 0.17 1.78 0.26 ;
  END
END DFFNRX4H7R

MACRO DFFNSRQX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNSRQX1H7R 0 0 ;
  SIZE 6.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.4 1.48 ;
        RECT 5.85 1.05 5.94 1.48 ;
        RECT 5.055 1.24 5.195 1.48 ;
        RECT 4.215 1.24 4.355 1.48 ;
        RECT 1.425 1.24 1.565 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.4 0.08 ;
        RECT 5.755 -0.08 5.895 0.305 ;
        RECT 4.96 -0.08 5.1 0.175 ;
        RECT 1.42 -0.08 1.56 0.175 ;
        RECT 0.36 -0.08 0.5 0.175 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.595 0.35 0.825 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.455 0.62 0.66 ;
        RECT 0.425 0.455 0.62 0.545 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.135 1.03 6.345 1.12 ;
        RECT 6.2 0.24 6.345 1.12 ;
        RECT 6.07 0.24 6.345 0.33 ;
        RECT 6.07 0.19 6.16 0.33 ;
      LAYER MET2 ;
        RECT 6.25 0.425 6.35 0.96 ;
      LAYER VIA1 ;
        RECT 6.255 0.655 6.345 0.745 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.82 0.45 4.99 0.67 ;
      LAYER MET2 ;
        RECT 4.85 0.23 4.95 0.76 ;
      LAYER VIA1 ;
        RECT 4.855 0.455 4.945 0.545 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.17 0.555 5.38 0.79 ;
      LAYER MET2 ;
        RECT 5.25 0.425 5.35 0.96 ;
      LAYER VIA1 ;
        RECT 5.255 0.655 5.345 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 4.473 1.14 4.934 1.23 ;
      RECT 3.765 1.14 4.095 1.23 ;
      RECT 4.431 1.14 4.976 1.209 ;
      RECT 3.765 1.14 4.137 1.209 ;
      RECT 4.393 1.14 5.014 1.169 ;
      RECT 3.765 1.14 4.175 1.169 ;
      RECT 5.67 0.855 5.76 1.15 ;
      RECT 4.896 1.121 5.76 1.15 ;
      RECT 4.976 1.06 5.76 1.15 ;
      RECT 4.057 1.121 4.511 1.15 ;
      RECT 4.934 1.081 5.76 1.15 ;
      RECT 4.095 1.081 4.473 1.15 ;
      RECT 4.137 1.06 4.431 1.15 ;
      RECT 5.67 0.855 6.005 0.945 ;
      RECT 5.915 0.405 6.005 0.945 ;
      RECT 5.915 0.56 6.09 0.7 ;
      RECT 5.53 0.405 6.005 0.495 ;
      RECT 5.53 0.22 5.62 0.495 ;
      RECT 4.55 0.96 4.858 1.05 ;
      RECT 4.508 0.96 4.9 1.029 ;
      RECT 4.47 0.96 4.938 0.989 ;
      RECT 5.475 0.585 5.565 0.97 ;
      RECT 3.285 0.71 3.375 0.97 ;
      RECT 4.82 0.941 5.565 0.97 ;
      RECT 4.9 0.88 5.565 0.97 ;
      RECT 4.165 0.941 4.588 0.97 ;
      RECT 4.858 0.901 5.565 0.97 ;
      RECT 4.165 0.901 4.55 0.97 ;
      RECT 4.165 0.88 4.508 0.97 ;
      RECT 4.165 0.71 4.255 0.97 ;
      RECT 3.285 0.71 4.255 0.8 ;
      RECT 3.82 0.35 3.91 0.8 ;
      RECT 5.475 0.585 5.825 0.675 ;
      RECT 3.105 0.35 4.47 0.44 ;
      RECT 4.863 0.265 5.39 0.355 ;
      RECT 5.3 0.205 5.39 0.355 ;
      RECT 4.852 0.221 4.863 0.35 ;
      RECT 2.23 0.17 2.32 0.345 ;
      RECT 4.806 0.193 4.852 0.321 ;
      RECT 4.768 0.246 4.901 0.279 ;
      RECT 2.23 0.17 4.806 0.26 ;
      RECT 4.64 0.78 4.78 0.87 ;
      RECT 4.64 0.35 4.73 0.87 ;
      RECT 4.12 0.53 4.73 0.62 ;
      RECT 4.59 0.35 4.73 0.62 ;
      RECT 2.155 1.14 3.555 1.23 ;
      RECT 3.465 0.89 3.555 1.23 ;
      RECT 3.465 0.89 4.075 0.98 ;
      RECT 1.941 0.96 3.195 1.05 ;
      RECT 3.105 0.53 3.195 1.05 ;
      RECT 1.899 0.901 1.941 1.029 ;
      RECT 1.871 0.96 3.195 0.994 ;
      RECT 1.755 0.96 3.195 0.98 ;
      RECT 1.04 0.88 1.899 0.97 ;
      RECT 1.04 0.941 1.979 0.97 ;
      RECT 1.04 0.538 1.13 0.97 ;
      RECT 3.105 0.53 3.73 0.62 ;
      RECT 1.04 0.538 1.156 0.586 ;
      RECT 1.086 0.493 1.194 0.554 ;
      RECT 1.086 0.493 1.713 0.535 ;
      RECT 1.13 0.458 1.759 0.512 ;
      RECT 1.156 0.445 1.808 0.459 ;
      RECT 1.759 0.355 1.77 0.484 ;
      RECT 1.675 0.426 1.808 0.459 ;
      RECT 1.713 0.384 1.759 0.512 ;
      RECT 1.77 0.35 1.91 0.44 ;
      RECT 2.018 0.78 3.015 0.87 ;
      RECT 2.925 0.35 3.015 0.87 ;
      RECT 1.976 0.721 2.018 0.849 ;
      RECT 1.938 0.78 3.015 0.809 ;
      RECT 1.275 0.7 1.976 0.79 ;
      RECT 1.275 0.761 2.056 0.79 ;
      RECT 2.485 0.35 3.015 0.44 ;
      RECT 0.045 0.915 0.16 1.16 ;
      RECT 0.045 0.915 0.77 1.005 ;
      RECT 0.68 0.74 0.77 1.005 ;
      RECT 0.045 0.24 0.135 1.16 ;
      RECT 2.126 0.53 2.835 0.62 ;
      RECT 2.09 0.474 2.126 0.602 ;
      RECT 2.046 0.511 2.164 0.562 ;
      RECT 2 0.17 2.09 0.517 ;
      RECT 1.344 0.265 1.637 0.355 ;
      RECT 0.045 0.265 0.68 0.355 ;
      RECT 0.59 0.17 0.68 0.355 ;
      RECT 1.333 0.221 1.344 0.35 ;
      RECT 1.333 0.265 1.683 0.332 ;
      RECT 1.287 0.193 1.333 0.321 ;
      RECT 1.599 0.246 1.732 0.279 ;
      RECT 1.683 0.175 1.694 0.304 ;
      RECT 1.249 0.246 1.382 0.279 ;
      RECT 0.045 0.24 0.195 0.355 ;
      RECT 1.694 0.17 2.09 0.26 ;
      RECT 0.59 0.17 1.287 0.26 ;
      RECT 1.637 0.204 2.09 0.26 ;
      RECT 1.683 1.14 2.065 1.23 ;
      RECT 1.641 1.081 1.683 1.209 ;
      RECT 0.755 1.095 0.95 1.185 ;
      RECT 0.86 0.35 0.95 1.185 ;
      RECT 1.603 1.14 2.065 1.169 ;
      RECT 0.86 1.06 1.641 1.15 ;
      RECT 0.755 1.121 1.721 1.15 ;
      RECT 0.86 0.35 1.005 0.44 ;
  END
END DFFNSRQX1H7R

MACRO DFFNSRQX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNSRQX2H7R 0 0 ;
  SIZE 6.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.6 1.48 ;
        RECT 6.42 1.005 6.51 1.48 ;
        RECT 5.85 1.05 5.94 1.48 ;
        RECT 5.055 1.24 5.195 1.48 ;
        RECT 4.215 1.24 4.355 1.48 ;
        RECT 1.425 1.24 1.565 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.6 0.08 ;
        RECT 6.38 -0.08 6.47 0.33 ;
        RECT 5.755 -0.08 5.895 0.305 ;
        RECT 4.96 -0.08 5.1 0.175 ;
        RECT 1.42 -0.08 1.56 0.175 ;
        RECT 0.36 -0.08 0.5 0.175 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.6 0.35 0.795 ;
        RECT 0.225 0.565 0.315 0.795 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.445 0.62 0.66 ;
        RECT 0.425 0.445 0.62 0.55 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.2 0.53 6.345 0.805 ;
        RECT 6.135 1.03 6.29 1.12 ;
        RECT 6.2 0.24 6.29 1.12 ;
        RECT 6.07 0.24 6.29 0.33 ;
        RECT 6.07 0.19 6.16 0.33 ;
      LAYER MET2 ;
        RECT 6.25 0.425 6.35 0.96 ;
      LAYER VIA1 ;
        RECT 6.255 0.655 6.345 0.745 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.82 0.45 4.99 0.67 ;
      LAYER MET2 ;
        RECT 4.85 0.23 4.95 0.76 ;
      LAYER VIA1 ;
        RECT 4.855 0.455 4.945 0.545 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.17 0.555 5.38 0.79 ;
      LAYER MET2 ;
        RECT 5.25 0.425 5.35 0.96 ;
      LAYER VIA1 ;
        RECT 5.255 0.655 5.345 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 4.473 1.14 4.934 1.23 ;
      RECT 3.765 1.14 4.095 1.23 ;
      RECT 4.431 1.14 4.976 1.209 ;
      RECT 3.765 1.14 4.137 1.209 ;
      RECT 4.393 1.14 5.014 1.169 ;
      RECT 3.765 1.14 4.175 1.169 ;
      RECT 5.67 0.855 5.76 1.15 ;
      RECT 4.896 1.121 5.76 1.15 ;
      RECT 4.976 1.06 5.76 1.15 ;
      RECT 4.057 1.121 4.511 1.15 ;
      RECT 4.934 1.081 5.76 1.15 ;
      RECT 4.095 1.081 4.473 1.15 ;
      RECT 4.137 1.06 4.431 1.15 ;
      RECT 5.67 0.855 6.005 0.945 ;
      RECT 5.915 0.405 6.005 0.945 ;
      RECT 5.915 0.56 6.09 0.7 ;
      RECT 5.53 0.405 6.005 0.495 ;
      RECT 5.53 0.22 5.62 0.495 ;
      RECT 4.55 0.96 4.858 1.05 ;
      RECT 4.508 0.96 4.9 1.029 ;
      RECT 4.47 0.96 4.938 0.989 ;
      RECT 5.475 0.585 5.565 0.97 ;
      RECT 3.285 0.71 3.375 0.97 ;
      RECT 4.82 0.941 5.565 0.97 ;
      RECT 4.9 0.88 5.565 0.97 ;
      RECT 4.165 0.941 4.588 0.97 ;
      RECT 4.858 0.901 5.565 0.97 ;
      RECT 4.165 0.901 4.55 0.97 ;
      RECT 4.165 0.88 4.508 0.97 ;
      RECT 4.165 0.71 4.255 0.97 ;
      RECT 3.285 0.71 4.255 0.8 ;
      RECT 3.82 0.35 3.91 0.8 ;
      RECT 5.475 0.585 5.825 0.675 ;
      RECT 3.105 0.35 4.47 0.44 ;
      RECT 4.863 0.265 5.39 0.355 ;
      RECT 5.3 0.205 5.39 0.355 ;
      RECT 4.852 0.221 4.863 0.35 ;
      RECT 2.23 0.17 2.32 0.345 ;
      RECT 4.806 0.193 4.852 0.321 ;
      RECT 4.768 0.246 4.901 0.279 ;
      RECT 2.23 0.17 4.806 0.26 ;
      RECT 4.64 0.78 4.78 0.87 ;
      RECT 4.64 0.35 4.73 0.87 ;
      RECT 4.12 0.53 4.73 0.62 ;
      RECT 4.59 0.35 4.73 0.62 ;
      RECT 2.155 1.14 3.555 1.23 ;
      RECT 3.465 0.89 3.555 1.23 ;
      RECT 3.465 0.89 4.075 0.98 ;
      RECT 1.941 0.96 3.195 1.05 ;
      RECT 3.105 0.53 3.195 1.05 ;
      RECT 1.899 0.901 1.941 1.029 ;
      RECT 1.871 0.96 3.195 0.994 ;
      RECT 1.755 0.96 3.195 0.98 ;
      RECT 1.04 0.88 1.899 0.97 ;
      RECT 1.04 0.941 1.979 0.97 ;
      RECT 1.04 0.538 1.13 0.97 ;
      RECT 3.105 0.53 3.73 0.62 ;
      RECT 1.04 0.538 1.156 0.586 ;
      RECT 1.086 0.493 1.194 0.554 ;
      RECT 1.086 0.493 1.713 0.535 ;
      RECT 1.13 0.458 1.759 0.512 ;
      RECT 1.156 0.445 1.808 0.459 ;
      RECT 1.759 0.355 1.77 0.484 ;
      RECT 1.675 0.426 1.808 0.459 ;
      RECT 1.713 0.384 1.759 0.512 ;
      RECT 1.77 0.35 1.91 0.44 ;
      RECT 2.018 0.78 3.015 0.87 ;
      RECT 2.925 0.35 3.015 0.87 ;
      RECT 1.976 0.721 2.018 0.849 ;
      RECT 1.938 0.78 3.015 0.809 ;
      RECT 1.275 0.7 1.976 0.79 ;
      RECT 1.275 0.761 2.056 0.79 ;
      RECT 2.485 0.35 3.015 0.44 ;
      RECT 0.045 0.915 0.16 1.16 ;
      RECT 0.045 0.915 0.77 1.005 ;
      RECT 0.68 0.74 0.77 1.005 ;
      RECT 0.045 0.24 0.135 1.16 ;
      RECT 2.126 0.53 2.835 0.62 ;
      RECT 2.09 0.474 2.126 0.602 ;
      RECT 2.046 0.511 2.164 0.562 ;
      RECT 2 0.17 2.09 0.517 ;
      RECT 1.344 0.265 1.637 0.355 ;
      RECT 0.045 0.265 0.68 0.355 ;
      RECT 0.59 0.17 0.68 0.355 ;
      RECT 1.333 0.221 1.344 0.35 ;
      RECT 1.333 0.265 1.683 0.332 ;
      RECT 1.287 0.193 1.333 0.321 ;
      RECT 1.599 0.246 1.732 0.279 ;
      RECT 1.683 0.175 1.694 0.304 ;
      RECT 1.249 0.246 1.382 0.279 ;
      RECT 0.045 0.24 0.195 0.355 ;
      RECT 1.694 0.17 2.09 0.26 ;
      RECT 0.59 0.17 1.287 0.26 ;
      RECT 1.637 0.204 2.09 0.26 ;
      RECT 1.683 1.14 2.065 1.23 ;
      RECT 1.641 1.081 1.683 1.209 ;
      RECT 0.755 1.095 0.95 1.185 ;
      RECT 0.86 0.35 0.95 1.185 ;
      RECT 1.603 1.14 2.065 1.169 ;
      RECT 0.86 1.06 1.641 1.15 ;
      RECT 0.755 1.121 1.721 1.15 ;
      RECT 0.86 0.35 1.005 0.44 ;
  END
END DFFNSRQX2H7R

MACRO DFFNSRX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNSRX0P5H7R 0 0 ;
  SIZE 7.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7.2 1.48 ;
        RECT 7.02 1.04 7.11 1.48 ;
        RECT 6.465 1.24 6.605 1.48 ;
        RECT 5.85 1.05 5.94 1.48 ;
        RECT 5.055 1.24 5.195 1.48 ;
        RECT 4.215 1.24 4.355 1.48 ;
        RECT 1.425 1.24 1.565 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7.2 0.08 ;
        RECT 6.39 -0.08 6.48 0.33 ;
        RECT 5.755 -0.08 5.895 0.305 ;
        RECT 4.96 -0.08 5.1 0.175 ;
        RECT 1.42 -0.08 1.56 0.175 ;
        RECT 0.36 -0.08 0.5 0.175 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.6 0.35 0.795 ;
        RECT 0.225 0.51 0.315 0.795 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.445 0.62 0.66 ;
        RECT 0.425 0.445 0.62 0.55 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.77 0.34 6.86 1.18 ;
        RECT 6.64 0.34 6.86 0.43 ;
        RECT 6.64 0.19 6.745 0.43 ;
      LAYER MET2 ;
        RECT 6.65 0.18 6.75 0.56 ;
      LAYER VIA1 ;
        RECT 6.655 0.255 6.745 0.345 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.195 0.625 6.35 0.92 ;
        RECT 6.095 0.625 6.35 0.765 ;
        RECT 6.095 0.215 6.185 0.765 ;
        RECT 6.005 0.215 6.185 0.305 ;
      LAYER MET2 ;
        RECT 6.25 0.425 6.35 0.96 ;
      LAYER VIA1 ;
        RECT 6.255 0.655 6.345 0.745 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.82 0.45 4.99 0.67 ;
      LAYER MET2 ;
        RECT 4.85 0.23 4.95 0.76 ;
      LAYER VIA1 ;
        RECT 4.855 0.455 4.945 0.545 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.17 0.555 5.38 0.79 ;
      LAYER MET2 ;
        RECT 5.25 0.425 5.35 0.96 ;
      LAYER VIA1 ;
        RECT 5.255 0.655 5.345 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 4.473 1.14 4.934 1.23 ;
      RECT 3.765 1.14 4.095 1.23 ;
      RECT 4.431 1.14 4.976 1.209 ;
      RECT 3.765 1.14 4.137 1.209 ;
      RECT 4.393 1.14 5.014 1.169 ;
      RECT 3.765 1.14 4.175 1.169 ;
      RECT 5.67 0.855 5.76 1.15 ;
      RECT 4.896 1.121 5.76 1.15 ;
      RECT 4.976 1.06 5.76 1.15 ;
      RECT 4.057 1.121 4.511 1.15 ;
      RECT 4.934 1.081 5.76 1.15 ;
      RECT 4.095 1.081 4.473 1.15 ;
      RECT 6.118 1.01 6.66 1.1 ;
      RECT 6.57 0.56 6.66 1.1 ;
      RECT 6.097 0.961 6.118 1.09 ;
      RECT 4.137 1.06 4.431 1.15 ;
      RECT 6.051 0.928 6.097 1.056 ;
      RECT 6.005 0.882 6.051 1.01 ;
      RECT 6.005 0.991 6.156 1.01 ;
      RECT 5.963 0.405 6.005 0.966 ;
      RECT 5.915 0.405 6.005 0.945 ;
      RECT 5.67 0.855 6.005 0.945 ;
      RECT 5.53 0.405 6.005 0.495 ;
      RECT 5.53 0.24 5.62 0.495 ;
      RECT 4.55 0.96 4.858 1.05 ;
      RECT 4.508 0.96 4.9 1.029 ;
      RECT 4.47 0.96 4.938 0.989 ;
      RECT 5.475 0.585 5.565 0.97 ;
      RECT 3.285 0.71 3.375 0.97 ;
      RECT 4.82 0.941 5.565 0.97 ;
      RECT 4.9 0.88 5.565 0.97 ;
      RECT 4.165 0.941 4.588 0.97 ;
      RECT 4.858 0.901 5.565 0.97 ;
      RECT 4.165 0.901 4.55 0.97 ;
      RECT 4.165 0.88 4.508 0.97 ;
      RECT 4.165 0.71 4.255 0.97 ;
      RECT 3.285 0.71 4.255 0.8 ;
      RECT 3.82 0.35 3.91 0.8 ;
      RECT 5.475 0.585 5.825 0.675 ;
      RECT 3.105 0.35 4.47 0.44 ;
      RECT 4.863 0.265 5.415 0.355 ;
      RECT 4.852 0.221 4.863 0.35 ;
      RECT 2.23 0.17 2.32 0.345 ;
      RECT 4.806 0.193 4.852 0.321 ;
      RECT 4.768 0.246 4.901 0.279 ;
      RECT 2.23 0.17 4.806 0.26 ;
      RECT 4.64 0.78 4.78 0.87 ;
      RECT 4.64 0.35 4.73 0.87 ;
      RECT 4.12 0.53 4.73 0.62 ;
      RECT 4.59 0.35 4.73 0.62 ;
      RECT 2.155 1.14 3.555 1.23 ;
      RECT 3.465 0.89 3.555 1.23 ;
      RECT 3.465 0.89 4.075 0.98 ;
      RECT 1.941 0.96 3.195 1.05 ;
      RECT 3.105 0.53 3.195 1.05 ;
      RECT 1.899 0.901 1.941 1.029 ;
      RECT 1.871 0.96 3.195 0.994 ;
      RECT 1.755 0.96 3.195 0.98 ;
      RECT 1.04 0.88 1.899 0.97 ;
      RECT 1.04 0.941 1.979 0.97 ;
      RECT 1.04 0.538 1.13 0.97 ;
      RECT 3.105 0.53 3.73 0.62 ;
      RECT 1.04 0.538 1.156 0.586 ;
      RECT 1.086 0.493 1.194 0.554 ;
      RECT 1.086 0.493 1.713 0.535 ;
      RECT 1.13 0.458 1.759 0.512 ;
      RECT 1.156 0.445 1.808 0.459 ;
      RECT 1.759 0.355 1.77 0.484 ;
      RECT 1.675 0.426 1.808 0.459 ;
      RECT 1.713 0.384 1.759 0.512 ;
      RECT 1.77 0.35 1.91 0.44 ;
      RECT 2.018 0.78 3.015 0.87 ;
      RECT 2.925 0.35 3.015 0.87 ;
      RECT 1.976 0.721 2.018 0.849 ;
      RECT 1.938 0.78 3.015 0.809 ;
      RECT 1.275 0.7 1.976 0.79 ;
      RECT 1.275 0.761 2.056 0.79 ;
      RECT 2.485 0.35 3.015 0.44 ;
      RECT 0.045 0.915 0.16 1.105 ;
      RECT 0.045 0.915 0.77 1.005 ;
      RECT 0.68 0.74 0.77 1.005 ;
      RECT 0.045 0.265 0.135 1.105 ;
      RECT 2.126 0.53 2.835 0.62 ;
      RECT 2.09 0.474 2.126 0.602 ;
      RECT 2.046 0.511 2.164 0.562 ;
      RECT 2 0.17 2.09 0.517 ;
      RECT 1.344 0.265 1.637 0.355 ;
      RECT 0.045 0.265 0.68 0.355 ;
      RECT 0.59 0.17 0.68 0.355 ;
      RECT 1.333 0.221 1.344 0.35 ;
      RECT 1.333 0.265 1.683 0.332 ;
      RECT 1.287 0.193 1.333 0.321 ;
      RECT 1.599 0.246 1.732 0.279 ;
      RECT 1.683 0.175 1.694 0.304 ;
      RECT 1.249 0.246 1.382 0.279 ;
      RECT 1.694 0.17 2.09 0.26 ;
      RECT 0.59 0.17 1.287 0.26 ;
      RECT 1.637 0.204 2.09 0.26 ;
      RECT 1.683 1.14 2.065 1.23 ;
      RECT 1.641 1.081 1.683 1.209 ;
      RECT 0.755 1.095 0.95 1.185 ;
      RECT 0.86 0.35 0.95 1.185 ;
      RECT 1.603 1.14 2.065 1.169 ;
      RECT 0.86 1.06 1.641 1.15 ;
      RECT 0.755 1.121 1.721 1.15 ;
      RECT 0.86 0.35 1.005 0.44 ;
  END
END DFFNSRX0P5H7R

MACRO DFFNSRX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNSRX1H7R 0 0 ;
  SIZE 7.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7.2 1.48 ;
        RECT 7.02 1.005 7.11 1.48 ;
        RECT 6.465 1.24 6.605 1.48 ;
        RECT 5.85 1.05 5.94 1.48 ;
        RECT 5.055 1.24 5.195 1.48 ;
        RECT 4.215 1.24 4.355 1.48 ;
        RECT 1.425 1.24 1.565 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7.2 0.08 ;
        RECT 6.95 -0.08 7.04 0.33 ;
        RECT 6.28 -0.08 6.37 0.33 ;
        RECT 5.755 -0.08 5.895 0.305 ;
        RECT 4.96 -0.08 5.1 0.175 ;
        RECT 1.42 -0.08 1.56 0.175 ;
        RECT 0.36 -0.08 0.5 0.175 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.6 0.35 0.795 ;
        RECT 0.225 0.51 0.315 0.795 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.445 0.62 0.66 ;
        RECT 0.425 0.445 0.62 0.55 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.77 0.34 6.86 1.145 ;
        RECT 6.64 0.34 6.86 0.43 ;
        RECT 6.64 0.19 6.745 0.43 ;
      LAYER MET2 ;
        RECT 6.65 0.18 6.75 0.56 ;
      LAYER VIA1 ;
        RECT 6.655 0.255 6.745 0.345 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.195 0.625 6.35 0.92 ;
        RECT 6.095 0.625 6.35 0.765 ;
        RECT 6.095 0.215 6.185 0.765 ;
        RECT 6.005 0.215 6.185 0.305 ;
      LAYER MET2 ;
        RECT 6.25 0.425 6.35 0.96 ;
      LAYER VIA1 ;
        RECT 6.255 0.655 6.345 0.745 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.82 0.455 4.99 0.67 ;
      LAYER MET2 ;
        RECT 4.85 0.23 4.95 0.76 ;
      LAYER VIA1 ;
        RECT 4.855 0.455 4.945 0.545 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.17 0.555 5.38 0.79 ;
      LAYER MET2 ;
        RECT 5.25 0.425 5.35 0.96 ;
      LAYER VIA1 ;
        RECT 5.255 0.655 5.345 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 4.473 1.14 4.934 1.23 ;
      RECT 3.765 1.14 4.095 1.23 ;
      RECT 4.431 1.14 4.976 1.209 ;
      RECT 3.765 1.14 4.137 1.209 ;
      RECT 4.393 1.14 5.014 1.169 ;
      RECT 3.765 1.14 4.175 1.169 ;
      RECT 5.67 0.855 5.76 1.15 ;
      RECT 4.896 1.121 5.76 1.15 ;
      RECT 4.976 1.06 5.76 1.15 ;
      RECT 4.057 1.121 4.511 1.15 ;
      RECT 4.934 1.081 5.76 1.15 ;
      RECT 4.095 1.081 4.473 1.15 ;
      RECT 6.118 1.01 6.66 1.1 ;
      RECT 6.57 0.56 6.66 1.1 ;
      RECT 6.097 0.961 6.118 1.09 ;
      RECT 4.137 1.06 4.431 1.15 ;
      RECT 6.051 0.928 6.097 1.056 ;
      RECT 6.005 0.882 6.051 1.01 ;
      RECT 6.005 0.991 6.156 1.01 ;
      RECT 5.963 0.405 6.005 0.966 ;
      RECT 5.915 0.405 6.005 0.945 ;
      RECT 5.67 0.855 6.005 0.945 ;
      RECT 5.53 0.405 6.005 0.495 ;
      RECT 5.53 0.24 5.62 0.495 ;
      RECT 4.55 0.96 4.858 1.05 ;
      RECT 4.508 0.96 4.9 1.029 ;
      RECT 4.47 0.96 4.938 0.989 ;
      RECT 5.475 0.585 5.565 0.97 ;
      RECT 3.285 0.71 3.375 0.97 ;
      RECT 4.82 0.941 5.565 0.97 ;
      RECT 4.9 0.88 5.565 0.97 ;
      RECT 4.165 0.941 4.588 0.97 ;
      RECT 4.858 0.901 5.565 0.97 ;
      RECT 4.165 0.901 4.55 0.97 ;
      RECT 4.165 0.88 4.508 0.97 ;
      RECT 4.165 0.71 4.255 0.97 ;
      RECT 3.285 0.71 4.255 0.8 ;
      RECT 3.82 0.35 3.91 0.8 ;
      RECT 5.475 0.585 5.825 0.675 ;
      RECT 3.105 0.35 4.47 0.44 ;
      RECT 4.863 0.265 5.415 0.355 ;
      RECT 4.852 0.221 4.863 0.35 ;
      RECT 2.23 0.17 2.32 0.345 ;
      RECT 4.806 0.193 4.852 0.321 ;
      RECT 4.768 0.246 4.901 0.279 ;
      RECT 2.23 0.17 4.806 0.26 ;
      RECT 4.64 0.78 4.78 0.87 ;
      RECT 4.64 0.35 4.73 0.87 ;
      RECT 4.12 0.53 4.73 0.62 ;
      RECT 4.59 0.35 4.73 0.62 ;
      RECT 2.155 1.14 3.555 1.23 ;
      RECT 3.465 0.89 3.555 1.23 ;
      RECT 3.465 0.89 4.075 0.98 ;
      RECT 1.941 0.96 3.195 1.05 ;
      RECT 3.105 0.53 3.195 1.05 ;
      RECT 1.899 0.901 1.941 1.029 ;
      RECT 1.871 0.96 3.195 0.994 ;
      RECT 1.755 0.96 3.195 0.98 ;
      RECT 1.04 0.88 1.899 0.97 ;
      RECT 1.04 0.941 1.979 0.97 ;
      RECT 1.04 0.538 1.13 0.97 ;
      RECT 3.105 0.53 3.73 0.62 ;
      RECT 1.04 0.538 1.156 0.586 ;
      RECT 1.086 0.493 1.194 0.554 ;
      RECT 1.086 0.493 1.713 0.535 ;
      RECT 1.13 0.458 1.759 0.512 ;
      RECT 1.156 0.445 1.808 0.459 ;
      RECT 1.759 0.355 1.77 0.484 ;
      RECT 1.675 0.426 1.808 0.459 ;
      RECT 1.713 0.384 1.759 0.512 ;
      RECT 1.77 0.35 1.91 0.44 ;
      RECT 2.018 0.78 3.015 0.87 ;
      RECT 2.925 0.35 3.015 0.87 ;
      RECT 1.976 0.721 2.018 0.849 ;
      RECT 1.938 0.78 3.015 0.809 ;
      RECT 1.275 0.7 1.976 0.79 ;
      RECT 1.275 0.761 2.056 0.79 ;
      RECT 2.485 0.35 3.015 0.44 ;
      RECT 0.045 0.915 0.16 1.105 ;
      RECT 0.045 0.915 0.77 1.005 ;
      RECT 0.68 0.74 0.77 1.005 ;
      RECT 0.045 0.265 0.135 1.105 ;
      RECT 2.126 0.53 2.835 0.62 ;
      RECT 2.09 0.474 2.126 0.602 ;
      RECT 2.046 0.511 2.164 0.562 ;
      RECT 2 0.17 2.09 0.517 ;
      RECT 1.344 0.265 1.637 0.355 ;
      RECT 0.045 0.265 0.68 0.355 ;
      RECT 0.59 0.17 0.68 0.355 ;
      RECT 1.333 0.221 1.344 0.35 ;
      RECT 1.333 0.265 1.683 0.332 ;
      RECT 1.287 0.193 1.333 0.321 ;
      RECT 1.599 0.246 1.732 0.279 ;
      RECT 1.683 0.175 1.694 0.304 ;
      RECT 1.249 0.246 1.382 0.279 ;
      RECT 1.694 0.17 2.09 0.26 ;
      RECT 0.59 0.17 1.287 0.26 ;
      RECT 1.637 0.204 2.09 0.26 ;
      RECT 1.683 1.14 2.065 1.23 ;
      RECT 1.641 1.081 1.683 1.209 ;
      RECT 0.755 1.095 0.95 1.185 ;
      RECT 0.86 0.35 0.95 1.185 ;
      RECT 1.603 1.14 2.065 1.169 ;
      RECT 0.86 1.06 1.641 1.15 ;
      RECT 0.755 1.121 1.721 1.15 ;
      RECT 0.86 0.35 1.005 0.44 ;
  END
END DFFNSRX1H7R

MACRO DFFNSRX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNSRX2H7R 0 0 ;
  SIZE 7.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7.2 1.48 ;
        RECT 7.02 1.005 7.11 1.48 ;
        RECT 6.465 1.24 6.605 1.48 ;
        RECT 5.85 1.05 5.94 1.48 ;
        RECT 5.055 1.24 5.195 1.48 ;
        RECT 4.215 1.24 4.355 1.48 ;
        RECT 1.425 1.24 1.565 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7.2 0.08 ;
        RECT 6.95 -0.08 7.04 0.33 ;
        RECT 6.28 -0.08 6.37 0.33 ;
        RECT 5.755 -0.08 5.895 0.305 ;
        RECT 4.96 -0.08 5.1 0.175 ;
        RECT 1.42 -0.08 1.56 0.175 ;
        RECT 0.36 -0.08 0.5 0.175 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.595 0.35 0.825 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.455 0.62 0.66 ;
        RECT 0.425 0.455 0.62 0.545 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.77 0.34 6.86 1.145 ;
        RECT 6.64 0.34 6.86 0.43 ;
        RECT 6.64 0.19 6.745 0.43 ;
      LAYER MET2 ;
        RECT 6.65 0.18 6.75 0.56 ;
      LAYER VIA1 ;
        RECT 6.655 0.255 6.745 0.345 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.095 0.625 6.35 0.775 ;
        RECT 6.195 0.625 6.285 0.92 ;
        RECT 6.095 0.225 6.185 0.775 ;
        RECT 6.005 0.225 6.185 0.315 ;
      LAYER MET2 ;
        RECT 6.25 0.425 6.35 0.96 ;
      LAYER VIA1 ;
        RECT 6.255 0.655 6.345 0.745 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.82 0.455 4.99 0.67 ;
      LAYER MET2 ;
        RECT 4.85 0.23 4.95 0.76 ;
      LAYER VIA1 ;
        RECT 4.855 0.455 4.945 0.545 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.17 0.555 5.38 0.79 ;
      LAYER MET2 ;
        RECT 5.25 0.425 5.35 0.96 ;
      LAYER VIA1 ;
        RECT 5.255 0.655 5.345 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 4.473 1.14 4.934 1.23 ;
      RECT 3.765 1.14 4.095 1.23 ;
      RECT 4.431 1.14 4.976 1.209 ;
      RECT 3.765 1.14 4.137 1.209 ;
      RECT 4.393 1.14 5.014 1.169 ;
      RECT 3.765 1.14 4.175 1.169 ;
      RECT 5.67 0.855 5.76 1.15 ;
      RECT 4.896 1.121 5.76 1.15 ;
      RECT 4.976 1.06 5.76 1.15 ;
      RECT 4.057 1.121 4.511 1.15 ;
      RECT 4.934 1.081 5.76 1.15 ;
      RECT 4.095 1.081 4.473 1.15 ;
      RECT 6.118 1.01 6.66 1.1 ;
      RECT 6.57 0.56 6.66 1.1 ;
      RECT 6.097 0.961 6.118 1.09 ;
      RECT 4.137 1.06 4.431 1.15 ;
      RECT 6.051 0.928 6.097 1.056 ;
      RECT 6.005 0.882 6.051 1.01 ;
      RECT 6.005 0.991 6.156 1.01 ;
      RECT 5.963 0.405 6.005 0.966 ;
      RECT 5.915 0.405 6.005 0.945 ;
      RECT 5.67 0.855 6.005 0.945 ;
      RECT 5.53 0.405 6.005 0.495 ;
      RECT 5.53 0.24 5.62 0.495 ;
      RECT 4.55 0.96 4.858 1.05 ;
      RECT 4.508 0.96 4.9 1.029 ;
      RECT 4.47 0.96 4.938 0.989 ;
      RECT 5.475 0.585 5.565 0.97 ;
      RECT 3.285 0.71 3.375 0.97 ;
      RECT 4.82 0.941 5.565 0.97 ;
      RECT 4.9 0.88 5.565 0.97 ;
      RECT 4.165 0.941 4.588 0.97 ;
      RECT 4.858 0.901 5.565 0.97 ;
      RECT 4.165 0.901 4.55 0.97 ;
      RECT 4.165 0.88 4.508 0.97 ;
      RECT 4.165 0.71 4.255 0.97 ;
      RECT 3.285 0.71 4.255 0.8 ;
      RECT 3.82 0.35 3.91 0.8 ;
      RECT 5.475 0.585 5.825 0.675 ;
      RECT 3.105 0.35 4.47 0.44 ;
      RECT 4.863 0.265 5.415 0.355 ;
      RECT 4.852 0.221 4.863 0.35 ;
      RECT 2.23 0.17 2.32 0.345 ;
      RECT 4.806 0.193 4.852 0.321 ;
      RECT 4.768 0.246 4.901 0.279 ;
      RECT 2.23 0.17 4.806 0.26 ;
      RECT 4.64 0.78 4.78 0.87 ;
      RECT 4.64 0.35 4.73 0.87 ;
      RECT 4.12 0.53 4.73 0.62 ;
      RECT 4.59 0.35 4.73 0.62 ;
      RECT 2.155 1.14 3.555 1.23 ;
      RECT 3.465 0.89 3.555 1.23 ;
      RECT 3.465 0.89 4.075 0.98 ;
      RECT 1.941 0.96 3.195 1.05 ;
      RECT 3.105 0.53 3.195 1.05 ;
      RECT 1.899 0.901 1.941 1.029 ;
      RECT 1.871 0.96 3.195 0.994 ;
      RECT 1.755 0.96 3.195 0.98 ;
      RECT 1.04 0.88 1.899 0.97 ;
      RECT 1.04 0.941 1.979 0.97 ;
      RECT 1.04 0.538 1.13 0.97 ;
      RECT 3.105 0.53 3.73 0.62 ;
      RECT 1.04 0.538 1.156 0.586 ;
      RECT 1.086 0.493 1.194 0.554 ;
      RECT 1.086 0.493 1.713 0.535 ;
      RECT 1.13 0.458 1.759 0.512 ;
      RECT 1.156 0.445 1.808 0.459 ;
      RECT 1.759 0.355 1.77 0.484 ;
      RECT 1.675 0.426 1.808 0.459 ;
      RECT 1.713 0.384 1.759 0.512 ;
      RECT 1.77 0.35 1.91 0.44 ;
      RECT 2.018 0.78 3.015 0.87 ;
      RECT 2.925 0.35 3.015 0.87 ;
      RECT 1.976 0.721 2.018 0.849 ;
      RECT 1.938 0.78 3.015 0.809 ;
      RECT 1.275 0.7 1.976 0.79 ;
      RECT 1.275 0.761 2.056 0.79 ;
      RECT 2.485 0.35 3.015 0.44 ;
      RECT 0.045 0.915 0.77 1.005 ;
      RECT 0.68 0.74 0.77 1.005 ;
      RECT 0.045 0.265 0.135 1.005 ;
      RECT 2.126 0.53 2.835 0.62 ;
      RECT 2.09 0.474 2.126 0.602 ;
      RECT 2.046 0.511 2.164 0.562 ;
      RECT 2 0.17 2.09 0.517 ;
      RECT 1.344 0.265 1.637 0.355 ;
      RECT 0.045 0.265 0.68 0.355 ;
      RECT 0.59 0.17 0.68 0.355 ;
      RECT 1.333 0.221 1.344 0.35 ;
      RECT 1.333 0.265 1.683 0.332 ;
      RECT 1.287 0.193 1.333 0.321 ;
      RECT 1.599 0.246 1.732 0.279 ;
      RECT 1.683 0.175 1.694 0.304 ;
      RECT 1.249 0.246 1.382 0.279 ;
      RECT 1.694 0.17 2.09 0.26 ;
      RECT 0.59 0.17 1.287 0.26 ;
      RECT 1.637 0.204 2.09 0.26 ;
      RECT 1.683 1.14 2.065 1.23 ;
      RECT 1.641 1.081 1.683 1.209 ;
      RECT 0.755 1.095 0.95 1.185 ;
      RECT 0.86 0.35 0.95 1.185 ;
      RECT 1.603 1.14 2.065 1.169 ;
      RECT 0.86 1.06 1.641 1.15 ;
      RECT 0.755 1.121 1.721 1.15 ;
      RECT 0.86 0.35 1.005 0.44 ;
  END
END DFFNSRX2H7R

MACRO DFFNSX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNSX0P5H7R 0 0 ;
  SIZE 6.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.6 1.48 ;
        RECT 6.145 0.885 6.235 1.48 ;
        RECT 5.128 1.095 5.268 1.48 ;
        RECT 4.321 1.24 4.461 1.48 ;
        RECT 2.593 1.24 2.733 1.48 ;
        RECT 1.795 1.24 1.935 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.6 0.08 ;
        RECT 6.12 -0.08 6.26 0.32 ;
        RECT 5.128 -0.08 5.268 0.305 ;
        RECT 4.402 -0.08 4.542 0.305 ;
        RECT 1.825 -0.08 1.965 0.16 ;
        RECT 0.36 -0.08 0.5 0.175 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.47 0.405 0.825 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.52 0.625 0.745 0.778 ;
        RECT 0.52 0.475 0.61 0.778 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.872 0.215 5.977 0.945 ;
        RECT 5.8 0.215 5.977 0.405 ;
      LAYER MET2 ;
        RECT 5.85 0.18 5.95 0.56 ;
      LAYER VIA1 ;
        RECT 5.855 0.255 5.945 0.345 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.462 0.287 5.602 0.905 ;
        RECT 5.41 0.655 5.602 0.745 ;
      LAYER MET2 ;
        RECT 5.45 0.425 5.55 0.96 ;
      LAYER VIA1 ;
        RECT 5.455 0.655 5.545 0.745 ;
    END
  END QN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.334 0.638 4.576 0.798 ;
      LAYER MET2 ;
        RECT 4.45 0.425 4.55 0.96 ;
      LAYER VIA1 ;
        RECT 4.455 0.655 4.545 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 4.579 1.14 4.993 1.23 ;
      RECT 4.903 0.915 4.993 1.23 ;
      RECT 4.537 1.081 4.579 1.209 ;
      RECT 4.132 1.06 4.222 1.2 ;
      RECT 4.499 1.14 4.993 1.169 ;
      RECT 4.132 1.06 4.537 1.15 ;
      RECT 4.132 1.121 4.617 1.15 ;
      RECT 5.386 0.995 5.782 1.085 ;
      RECT 5.692 0.55 5.782 1.085 ;
      RECT 5.344 0.936 5.386 1.064 ;
      RECT 5.306 0.995 5.782 1.024 ;
      RECT 4.903 0.915 5.344 1.005 ;
      RECT 4.903 0.976 5.424 1.005 ;
      RECT 5.141 0.395 5.231 1.005 ;
      RECT 4.903 0.395 5.231 0.485 ;
      RECT 4.903 0.224 4.993 0.485 ;
      RECT 4.666 0.42 4.756 1.014 ;
      RECT 3.262 0.899 3.752 0.989 ;
      RECT 3.662 0.35 3.752 0.989 ;
      RECT 4.666 0.575 5.051 0.665 ;
      RECT 4.021 0.42 4.756 0.51 ;
      RECT 3.989 0.366 4.021 0.494 ;
      RECT 3.951 0.42 4.756 0.459 ;
      RECT 3.662 0.35 3.989 0.44 ;
      RECT 3.662 0.401 4.059 0.44 ;
      RECT 2.565 0.17 2.705 0.32 ;
      RECT 4.152 0.17 4.292 0.305 ;
      RECT 2.565 0.17 4.292 0.26 ;
      RECT 2.954 1.14 3.932 1.23 ;
      RECT 3.842 0.648 3.932 1.23 ;
      RECT 2.912 1.081 2.954 1.209 ;
      RECT 2.874 1.14 3.932 1.169 ;
      RECT 2.641 1.06 2.912 1.15 ;
      RECT 2.625 1.014 2.641 1.142 ;
      RECT 2.625 1.121 2.992 1.142 ;
      RECT 2.579 0.983 2.625 1.111 ;
      RECT 2.541 1.041 2.679 1.069 ;
      RECT 2.165 0.96 2.579 1.05 ;
      RECT 2.123 0.901 2.165 1.029 ;
      RECT 2.085 0.88 2.123 0.989 ;
      RECT 1.4 0.88 2.123 0.97 ;
      RECT 1.4 0.941 2.203 0.97 ;
      RECT 1.4 0.777 1.49 0.97 ;
      RECT 1.015 0.777 1.49 0.867 ;
      RECT 1.015 0.578 1.105 0.867 ;
      RECT 1.061 0.533 1.151 0.616 ;
      RECT 1.105 0.488 1.224 0.539 ;
      RECT 1.151 0.447 1.186 0.576 ;
      RECT 2.155 0.373 2.295 0.52 ;
      RECT 1.186 0.43 2.295 0.52 ;
      RECT 2.717 0.88 3.063 0.97 ;
      RECT 2.701 0.834 2.717 0.962 ;
      RECT 2.701 0.88 3.109 0.947 ;
      RECT 2.655 0.803 2.701 0.931 ;
      RECT 3.025 0.861 3.155 0.901 ;
      RECT 2.617 0.861 2.755 0.889 ;
      RECT 2.241 0.78 2.655 0.87 ;
      RECT 2.227 0.735 2.241 0.863 ;
      RECT 3.063 0.819 3.186 0.863 ;
      RECT 2.181 0.705 2.227 0.833 ;
      RECT 3.109 0.773 3.224 0.828 ;
      RECT 3.155 0.734 3.186 0.863 ;
      RECT 3.482 0.35 3.572 0.809 ;
      RECT 2.135 0.659 2.181 0.787 ;
      RECT 2.135 0.761 2.279 0.787 ;
      RECT 3.186 0.719 3.572 0.809 ;
      RECT 2.117 0.61 2.135 0.755 ;
      RECT 2.071 0.61 2.135 0.723 ;
      RECT 1.634 0.61 2.135 0.7 ;
      RECT 2.86 0.35 3.572 0.44 ;
      RECT 0.606 1.137 1.13 1.227 ;
      RECT 0.045 0.915 0.185 1.16 ;
      RECT 0.606 0.915 0.696 1.227 ;
      RECT 0.045 0.915 0.696 1.005 ;
      RECT 0.045 0.27 0.135 1.16 ;
      RECT 2.385 0.539 3.392 0.629 ;
      RECT 2.385 0.17 2.475 0.629 ;
      RECT 0.045 0.27 0.68 0.36 ;
      RECT 0.59 0.17 0.68 0.36 ;
      RECT 1.586 0.25 2.041 0.34 ;
      RECT 1.544 0.25 2.083 0.319 ;
      RECT 1.506 0.25 2.121 0.279 ;
      RECT 2.083 0.17 2.475 0.26 ;
      RECT 2.003 0.231 2.475 0.26 ;
      RECT 2.041 0.191 2.083 0.319 ;
      RECT 0.59 0.231 1.624 0.26 ;
      RECT 0.59 0.191 1.586 0.26 ;
      RECT 0.59 0.17 1.544 0.26 ;
      RECT 2.089 1.14 2.503 1.23 ;
      RECT 2.047 1.081 2.089 1.209 ;
      RECT 2.009 1.14 2.503 1.169 ;
      RECT 1.22 1.06 2.047 1.15 ;
      RECT 1.22 1.121 2.127 1.15 ;
      RECT 1.22 0.957 1.31 1.15 ;
      RECT 0.81 0.957 1.31 1.047 ;
      RECT 0.835 0.355 0.925 1.047 ;
      RECT 0.835 0.355 1.043 0.445 ;
  END
END DFFNSX0P5H7R

MACRO DFFNSX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNSX1H7R 0 0 ;
  SIZE 6.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.6 1.48 ;
        RECT 6.145 0.975 6.235 1.48 ;
        RECT 5.128 1.095 5.268 1.48 ;
        RECT 4.321 1.24 4.461 1.48 ;
        RECT 2.593 1.24 2.733 1.48 ;
        RECT 1.795 1.24 1.935 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.6 0.08 ;
        RECT 6.12 -0.08 6.26 0.32 ;
        RECT 5.128 -0.08 5.268 0.305 ;
        RECT 4.402 -0.08 4.542 0.305 ;
        RECT 1.825 -0.08 1.965 0.16 ;
        RECT 0.36 -0.08 0.5 0.175 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.47 0.405 0.825 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.52 0.625 0.745 0.783 ;
        RECT 0.52 0.475 0.61 0.783 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.872 0.225 5.982 0.945 ;
        RECT 5.82 0.225 5.982 0.425 ;
      LAYER MET2 ;
        RECT 5.85 0.18 5.95 0.56 ;
      LAYER VIA1 ;
        RECT 5.855 0.255 5.945 0.345 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.462 0.287 5.602 0.905 ;
        RECT 5.41 0.655 5.602 0.745 ;
      LAYER MET2 ;
        RECT 5.45 0.425 5.55 0.96 ;
      LAYER VIA1 ;
        RECT 5.455 0.655 5.545 0.745 ;
    END
  END QN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.334 0.638 4.576 0.798 ;
      LAYER MET2 ;
        RECT 4.45 0.425 4.55 0.96 ;
      LAYER VIA1 ;
        RECT 4.455 0.655 4.545 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 4.579 1.14 4.993 1.23 ;
      RECT 4.903 0.915 4.993 1.23 ;
      RECT 4.537 1.081 4.579 1.209 ;
      RECT 4.132 1.06 4.222 1.2 ;
      RECT 4.499 1.14 4.993 1.169 ;
      RECT 4.132 1.06 4.537 1.15 ;
      RECT 4.132 1.121 4.617 1.15 ;
      RECT 5.386 0.995 5.782 1.085 ;
      RECT 5.692 0.55 5.782 1.085 ;
      RECT 5.344 0.936 5.386 1.064 ;
      RECT 5.306 0.995 5.782 1.024 ;
      RECT 4.903 0.915 5.344 1.005 ;
      RECT 4.903 0.976 5.424 1.005 ;
      RECT 5.141 0.395 5.231 1.005 ;
      RECT 4.903 0.395 5.231 0.485 ;
      RECT 4.903 0.224 4.993 0.485 ;
      RECT 4.666 0.42 4.756 1.014 ;
      RECT 3.262 0.899 3.752 0.989 ;
      RECT 3.662 0.35 3.752 0.989 ;
      RECT 4.666 0.575 5.051 0.665 ;
      RECT 4.021 0.42 4.756 0.51 ;
      RECT 3.989 0.366 4.021 0.494 ;
      RECT 3.951 0.42 4.756 0.459 ;
      RECT 3.662 0.35 3.989 0.44 ;
      RECT 3.662 0.401 4.059 0.44 ;
      RECT 2.565 0.17 2.705 0.32 ;
      RECT 4.152 0.17 4.292 0.305 ;
      RECT 2.565 0.17 4.292 0.26 ;
      RECT 2.954 1.14 3.932 1.23 ;
      RECT 3.842 0.648 3.932 1.23 ;
      RECT 2.912 1.081 2.954 1.209 ;
      RECT 2.874 1.14 3.932 1.169 ;
      RECT 2.641 1.06 2.912 1.15 ;
      RECT 2.625 1.014 2.641 1.142 ;
      RECT 2.625 1.121 2.992 1.142 ;
      RECT 2.579 0.983 2.625 1.111 ;
      RECT 2.541 1.041 2.679 1.069 ;
      RECT 2.165 0.96 2.579 1.05 ;
      RECT 2.123 0.901 2.165 1.029 ;
      RECT 2.085 0.88 2.123 0.989 ;
      RECT 1.4 0.88 2.123 0.97 ;
      RECT 1.4 0.941 2.203 0.97 ;
      RECT 1.4 0.777 1.49 0.97 ;
      RECT 1.015 0.777 1.49 0.867 ;
      RECT 1.015 0.578 1.105 0.867 ;
      RECT 1.061 0.533 1.151 0.616 ;
      RECT 1.105 0.488 1.224 0.539 ;
      RECT 1.151 0.447 1.186 0.576 ;
      RECT 2.155 0.373 2.295 0.52 ;
      RECT 1.186 0.43 2.295 0.52 ;
      RECT 2.717 0.88 3.063 0.97 ;
      RECT 2.701 0.834 2.717 0.962 ;
      RECT 2.701 0.88 3.109 0.947 ;
      RECT 2.655 0.803 2.701 0.931 ;
      RECT 3.025 0.861 3.155 0.901 ;
      RECT 2.617 0.861 2.755 0.889 ;
      RECT 2.241 0.78 2.655 0.87 ;
      RECT 2.227 0.735 2.241 0.863 ;
      RECT 3.063 0.819 3.186 0.863 ;
      RECT 2.181 0.705 2.227 0.833 ;
      RECT 3.109 0.773 3.224 0.828 ;
      RECT 3.155 0.734 3.186 0.863 ;
      RECT 3.482 0.35 3.572 0.809 ;
      RECT 2.135 0.659 2.181 0.787 ;
      RECT 2.135 0.761 2.279 0.787 ;
      RECT 3.186 0.719 3.572 0.809 ;
      RECT 2.117 0.61 2.135 0.755 ;
      RECT 2.071 0.61 2.135 0.723 ;
      RECT 1.634 0.61 2.135 0.7 ;
      RECT 2.86 0.35 3.572 0.44 ;
      RECT 0.606 1.137 1.13 1.227 ;
      RECT 0.045 0.915 0.185 1.16 ;
      RECT 0.606 0.915 0.696 1.227 ;
      RECT 0.045 0.915 0.696 1.005 ;
      RECT 0.045 0.27 0.135 1.16 ;
      RECT 2.385 0.539 3.392 0.629 ;
      RECT 2.385 0.17 2.475 0.629 ;
      RECT 0.045 0.27 0.68 0.36 ;
      RECT 0.59 0.17 0.68 0.36 ;
      RECT 1.586 0.25 2.041 0.34 ;
      RECT 1.544 0.25 2.083 0.319 ;
      RECT 1.506 0.25 2.121 0.279 ;
      RECT 2.083 0.17 2.475 0.26 ;
      RECT 2.003 0.231 2.475 0.26 ;
      RECT 2.041 0.191 2.083 0.319 ;
      RECT 0.59 0.231 1.624 0.26 ;
      RECT 0.59 0.191 1.586 0.26 ;
      RECT 0.59 0.17 1.544 0.26 ;
      RECT 2.089 1.14 2.503 1.23 ;
      RECT 2.047 1.081 2.089 1.209 ;
      RECT 2.009 1.14 2.503 1.169 ;
      RECT 1.22 1.06 2.047 1.15 ;
      RECT 1.22 1.121 2.127 1.15 ;
      RECT 1.22 0.957 1.31 1.15 ;
      RECT 0.81 0.957 1.31 1.047 ;
      RECT 0.835 0.355 0.925 1.047 ;
      RECT 0.835 0.355 1.043 0.445 ;
  END
END DFFNSX1H7R

MACRO DFFNSX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNSX2H7R 0 0 ;
  SIZE 6.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.6 1.48 ;
        RECT 6.145 1.055 6.235 1.48 ;
        RECT 5.128 1.095 5.268 1.48 ;
        RECT 4.321 1.24 4.461 1.48 ;
        RECT 2.593 1.24 2.733 1.48 ;
        RECT 1.795 1.24 1.935 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.6 0.08 ;
        RECT 6.12 -0.08 6.26 0.32 ;
        RECT 5.128 -0.08 5.268 0.305 ;
        RECT 4.402 -0.08 4.542 0.305 ;
        RECT 1.825 -0.08 1.965 0.16 ;
        RECT 0.36 -0.08 0.5 0.175 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.445 0.405 0.825 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.52 0.625 0.745 0.775 ;
        RECT 0.52 0.445 0.61 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.872 0.225 5.975 1.145 ;
        RECT 5.82 0.225 5.975 0.345 ;
      LAYER MET2 ;
        RECT 5.85 0.18 5.95 0.56 ;
      LAYER VIA1 ;
        RECT 5.855 0.255 5.945 0.345 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.462 0.287 5.602 0.905 ;
        RECT 5.43 0.625 5.602 0.775 ;
      LAYER MET2 ;
        RECT 5.45 0.425 5.55 0.96 ;
      LAYER VIA1 ;
        RECT 5.455 0.655 5.545 0.745 ;
    END
  END QN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.334 0.638 4.576 0.798 ;
      LAYER MET2 ;
        RECT 4.45 0.425 4.55 0.96 ;
      LAYER VIA1 ;
        RECT 4.455 0.655 4.545 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 4.579 1.14 4.993 1.23 ;
      RECT 4.903 0.915 4.993 1.23 ;
      RECT 4.537 1.081 4.579 1.209 ;
      RECT 4.132 1.06 4.222 1.2 ;
      RECT 4.499 1.14 4.993 1.169 ;
      RECT 4.132 1.06 4.537 1.15 ;
      RECT 4.132 1.121 4.617 1.15 ;
      RECT 5.386 0.995 5.782 1.085 ;
      RECT 5.692 0.55 5.782 1.085 ;
      RECT 5.344 0.936 5.386 1.064 ;
      RECT 5.306 0.995 5.782 1.024 ;
      RECT 4.903 0.915 5.344 1.005 ;
      RECT 4.903 0.976 5.424 1.005 ;
      RECT 5.141 0.395 5.231 1.005 ;
      RECT 4.903 0.395 5.231 0.485 ;
      RECT 4.903 0.224 4.993 0.485 ;
      RECT 4.666 0.42 4.756 1.014 ;
      RECT 3.262 0.899 3.752 0.989 ;
      RECT 3.662 0.35 3.752 0.989 ;
      RECT 4.666 0.575 5.051 0.665 ;
      RECT 4.021 0.42 4.756 0.51 ;
      RECT 3.989 0.366 4.021 0.494 ;
      RECT 3.951 0.42 4.756 0.459 ;
      RECT 3.662 0.35 3.989 0.44 ;
      RECT 3.662 0.401 4.059 0.44 ;
      RECT 2.565 0.17 2.705 0.32 ;
      RECT 4.152 0.17 4.292 0.305 ;
      RECT 2.565 0.17 4.292 0.26 ;
      RECT 2.954 1.14 3.932 1.23 ;
      RECT 3.842 0.648 3.932 1.23 ;
      RECT 2.912 1.081 2.954 1.209 ;
      RECT 2.874 1.14 3.932 1.169 ;
      RECT 2.641 1.06 2.912 1.15 ;
      RECT 2.625 1.014 2.641 1.142 ;
      RECT 2.625 1.121 2.992 1.142 ;
      RECT 2.579 0.983 2.625 1.111 ;
      RECT 2.541 1.041 2.679 1.069 ;
      RECT 2.165 0.96 2.579 1.05 ;
      RECT 2.123 0.901 2.165 1.029 ;
      RECT 2.085 0.88 2.123 0.989 ;
      RECT 1.4 0.88 2.123 0.97 ;
      RECT 1.4 0.941 2.203 0.97 ;
      RECT 1.4 0.777 1.49 0.97 ;
      RECT 1.015 0.777 1.49 0.867 ;
      RECT 1.015 0.578 1.105 0.867 ;
      RECT 1.061 0.533 1.151 0.616 ;
      RECT 1.105 0.488 1.224 0.539 ;
      RECT 1.151 0.447 1.186 0.576 ;
      RECT 2.155 0.373 2.295 0.52 ;
      RECT 1.186 0.43 2.295 0.52 ;
      RECT 2.717 0.88 3.063 0.97 ;
      RECT 2.701 0.834 2.717 0.962 ;
      RECT 2.701 0.88 3.109 0.947 ;
      RECT 2.655 0.803 2.701 0.931 ;
      RECT 3.025 0.861 3.155 0.901 ;
      RECT 2.617 0.861 2.755 0.889 ;
      RECT 2.241 0.78 2.655 0.87 ;
      RECT 2.227 0.735 2.241 0.863 ;
      RECT 3.063 0.819 3.186 0.863 ;
      RECT 2.181 0.705 2.227 0.833 ;
      RECT 3.109 0.773 3.224 0.828 ;
      RECT 3.155 0.734 3.186 0.863 ;
      RECT 3.482 0.35 3.572 0.809 ;
      RECT 2.135 0.659 2.181 0.787 ;
      RECT 2.135 0.761 2.279 0.787 ;
      RECT 3.186 0.719 3.572 0.809 ;
      RECT 2.117 0.61 2.135 0.755 ;
      RECT 2.071 0.61 2.135 0.723 ;
      RECT 1.634 0.61 2.135 0.7 ;
      RECT 2.86 0.35 3.572 0.44 ;
      RECT 0.606 1.137 1.13 1.227 ;
      RECT 0.045 0.915 0.185 1.16 ;
      RECT 0.606 0.915 0.696 1.227 ;
      RECT 0.045 0.915 0.696 1.005 ;
      RECT 0.045 0.225 0.135 1.16 ;
      RECT 2.385 0.539 3.392 0.629 ;
      RECT 2.385 0.17 2.475 0.629 ;
      RECT 0.045 0.265 0.68 0.355 ;
      RECT 0.59 0.17 0.68 0.355 ;
      RECT 1.586 0.25 2.041 0.34 ;
      RECT 1.544 0.25 2.083 0.319 ;
      RECT 1.506 0.25 2.121 0.279 ;
      RECT 0.045 0.225 0.185 0.355 ;
      RECT 2.083 0.17 2.475 0.26 ;
      RECT 2.003 0.231 2.475 0.26 ;
      RECT 2.041 0.191 2.083 0.319 ;
      RECT 0.59 0.231 1.624 0.26 ;
      RECT 0.59 0.191 1.586 0.26 ;
      RECT 0.59 0.17 1.544 0.26 ;
      RECT 2.089 1.14 2.503 1.23 ;
      RECT 2.047 1.081 2.089 1.209 ;
      RECT 2.009 1.14 2.503 1.169 ;
      RECT 1.22 1.06 2.047 1.15 ;
      RECT 1.22 1.121 2.127 1.15 ;
      RECT 1.22 0.957 1.31 1.15 ;
      RECT 0.81 0.957 1.31 1.047 ;
      RECT 0.835 0.355 0.925 1.047 ;
      RECT 0.835 0.355 1.043 0.445 ;
  END
END DFFNSX2H7R

MACRO DFFNX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNX0P5H7R 0 0 ;
  SIZE 5 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5 1.48 ;
        RECT 4.482 1.225 4.622 1.48 ;
        RECT 3.642 1.225 3.782 1.48 ;
        RECT 2.287 1.095 2.427 1.48 ;
        RECT 1.47 1.225 1.61 1.48 ;
        RECT 0.31 1.15 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5 0.08 ;
        RECT 4.482 -0.08 4.622 0.36 ;
        RECT 3.592 -0.08 3.732 0.34 ;
        RECT 2.302 -0.08 2.442 0.175 ;
        RECT 1.455 -0.08 1.595 0.16 ;
        RECT 0.325 -0.08 0.465 0.16 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.605 0.355 0.865 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.455 0.626 0.6 ;
        RECT 0.425 0.455 0.626 0.545 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.772 0.31 4.862 0.987 ;
        RECT 4.625 0.455 4.862 0.545 ;
      LAYER MET2 ;
        RECT 4.65 0.225 4.75 0.76 ;
      LAYER VIA1 ;
        RECT 4.655 0.455 4.745 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.987 0.865 4.127 1.04 ;
        RECT 3.625 0.865 4.127 0.955 ;
        RECT 3.625 0.455 3.972 0.545 ;
        RECT 3.882 0.35 3.972 0.545 ;
        RECT 3.625 0.455 3.715 0.955 ;
      LAYER MET2 ;
        RECT 3.65 0.23 3.75 0.76 ;
      LAYER VIA1 ;
        RECT 3.655 0.455 3.745 0.545 ;
    END
  END QN
  OBS
    LAYER MET1 ;
      RECT 3.915 1.14 4.346 1.23 ;
      RECT 3.904 1.096 3.915 1.225 ;
      RECT 3.904 1.14 4.392 1.207 ;
      RECT 3.858 1.068 3.904 1.196 ;
      RECT 4.308 1.121 4.422 1.169 ;
      RECT 3.82 1.121 3.953 1.154 ;
      RECT 3.092 1.045 3.858 1.135 ;
      RECT 4.346 1.079 4.468 1.131 ;
      RECT 4.392 1.041 4.422 1.169 ;
      RECT 4.422 0.587 4.512 1.086 ;
      RECT 3.092 0.395 3.182 1.135 ;
      RECT 2.807 0.395 3.182 0.485 ;
      RECT 4.242 0.31 4.332 0.987 ;
      RECT 3.807 0.654 4.332 0.744 ;
      RECT 0.585 1.14 1.055 1.23 ;
      RECT 0.585 0.96 0.675 1.23 ;
      RECT 0.07 0.96 0.675 1.05 ;
      RECT 0.07 0.25 0.16 1.05 ;
      RECT 3.272 0.17 3.362 0.816 ;
      RECT 2.223 0.265 2.604 0.355 ;
      RECT 2.212 0.221 2.223 0.35 ;
      RECT 1.377 0.25 1.671 0.34 ;
      RECT 0.07 0.25 0.681 0.34 ;
      RECT 2.212 0.265 2.65 0.332 ;
      RECT 2.166 0.193 2.212 0.321 ;
      RECT 1.335 0.25 1.713 0.319 ;
      RECT 1.297 0.25 1.751 0.279 ;
      RECT 2.566 0.246 2.699 0.279 ;
      RECT 2.65 0.175 2.661 0.304 ;
      RECT 2.128 0.246 2.261 0.279 ;
      RECT 2.661 0.17 3.362 0.26 ;
      RECT 1.713 0.17 2.166 0.26 ;
      RECT 1.671 0.191 1.713 0.319 ;
      RECT 0.591 0.231 1.415 0.26 ;
      RECT 2.604 0.204 3.362 0.26 ;
      RECT 1.633 0.231 2.223 0.26 ;
      RECT 0.591 0.191 1.377 0.26 ;
      RECT 0.591 0.17 1.335 0.26 ;
      RECT 1.743 1.14 2.152 1.23 ;
      RECT 2.062 0.845 2.152 1.23 ;
      RECT 1.732 1.096 1.743 1.225 ;
      RECT 1.686 1.068 1.732 1.196 ;
      RECT 1.648 1.121 1.781 1.154 ;
      RECT 1.145 1.045 1.686 1.135 ;
      RECT 1.145 0.745 1.235 1.135 ;
      RECT 2.062 0.845 2.985 0.935 ;
      RECT 2.895 0.74 2.985 0.935 ;
      RECT 2.627 0.445 2.717 0.935 ;
      RECT 1.065 0.745 1.235 0.835 ;
      RECT 2.035 0.445 2.717 0.535 ;
      RECT 1.799 0.37 1.889 1.03 ;
      RECT 1.35 0.865 1.889 0.955 ;
      RECT 1.35 0.625 1.44 0.955 ;
      RECT 1.799 0.665 2.537 0.755 ;
      RECT 1.774 0.37 1.914 0.46 ;
      RECT 0.85 0.37 0.94 1.03 ;
      RECT 1.61 0.532 1.7 0.7 ;
      RECT 1.576 0.447 1.61 0.575 ;
      RECT 1.538 0.487 1.656 0.539 ;
      RECT 0.85 0.43 1.576 0.52 ;
      RECT 0.85 0.37 1.03 0.52 ;
  END
END DFFNX0P5H7R

MACRO DFFNX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNX1H7R 0 0 ;
  SIZE 5 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5 1.48 ;
        RECT 4.482 1.225 4.622 1.48 ;
        RECT 3.642 1.225 3.782 1.48 ;
        RECT 2.287 1.062 2.427 1.48 ;
        RECT 1.47 1.225 1.61 1.48 ;
        RECT 0.31 1.15 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5 0.08 ;
        RECT 4.355 -0.08 4.495 0.335 ;
        RECT 3.592 -0.08 3.732 0.34 ;
        RECT 2.302 -0.08 2.442 0.175 ;
        RECT 1.455 -0.08 1.595 0.16 ;
        RECT 0.325 -0.08 0.465 0.16 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.605 0.355 0.865 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.455 0.626 0.6 ;
        RECT 0.425 0.455 0.626 0.545 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.772 0.455 4.862 0.987 ;
        RECT 4.625 0.455 4.862 0.545 ;
        RECT 4.625 0.31 4.72 0.545 ;
      LAYER MET2 ;
        RECT 4.65 0.225 4.75 0.76 ;
      LAYER VIA1 ;
        RECT 4.655 0.455 4.745 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.987 0.865 4.127 1.04 ;
        RECT 3.625 0.865 4.127 0.955 ;
        RECT 3.625 0.455 3.972 0.545 ;
        RECT 3.882 0.35 3.972 0.545 ;
        RECT 3.625 0.455 3.715 0.955 ;
      LAYER MET2 ;
        RECT 3.65 0.23 3.75 0.76 ;
      LAYER VIA1 ;
        RECT 3.655 0.455 3.745 0.545 ;
    END
  END QN
  OBS
    LAYER MET1 ;
      RECT 3.915 1.14 4.346 1.23 ;
      RECT 3.904 1.096 3.915 1.225 ;
      RECT 3.904 1.14 4.392 1.207 ;
      RECT 3.858 1.068 3.904 1.196 ;
      RECT 4.308 1.121 4.422 1.169 ;
      RECT 3.82 1.121 3.953 1.154 ;
      RECT 3.092 1.045 3.858 1.135 ;
      RECT 4.346 1.079 4.468 1.131 ;
      RECT 4.392 1.041 4.422 1.169 ;
      RECT 4.422 0.587 4.512 1.086 ;
      RECT 3.092 0.395 3.182 1.135 ;
      RECT 2.807 0.395 3.182 0.485 ;
      RECT 4.242 0.654 4.332 0.987 ;
      RECT 3.807 0.654 4.332 0.744 ;
      RECT 4.115 0.31 4.205 0.744 ;
      RECT 0.585 1.14 1.055 1.23 ;
      RECT 0.585 0.96 0.675 1.23 ;
      RECT 0.07 0.96 0.675 1.05 ;
      RECT 0.07 0.25 0.16 1.05 ;
      RECT 3.272 0.17 3.362 0.816 ;
      RECT 2.223 0.265 2.599 0.355 ;
      RECT 2.212 0.221 2.223 0.35 ;
      RECT 1.377 0.25 1.671 0.34 ;
      RECT 0.07 0.25 0.681 0.34 ;
      RECT 2.212 0.265 2.645 0.332 ;
      RECT 2.166 0.193 2.212 0.321 ;
      RECT 1.335 0.25 1.713 0.319 ;
      RECT 1.297 0.25 1.751 0.279 ;
      RECT 2.561 0.246 2.694 0.279 ;
      RECT 2.645 0.175 2.656 0.304 ;
      RECT 2.128 0.246 2.261 0.279 ;
      RECT 2.656 0.17 3.362 0.26 ;
      RECT 1.713 0.17 2.166 0.26 ;
      RECT 1.671 0.191 1.713 0.319 ;
      RECT 0.591 0.231 1.415 0.26 ;
      RECT 2.599 0.204 3.362 0.26 ;
      RECT 1.633 0.231 2.223 0.26 ;
      RECT 0.591 0.191 1.377 0.26 ;
      RECT 0.591 0.17 1.335 0.26 ;
      RECT 1.743 1.14 2.152 1.23 ;
      RECT 2.062 0.845 2.152 1.23 ;
      RECT 1.732 1.096 1.743 1.225 ;
      RECT 1.686 1.068 1.732 1.196 ;
      RECT 1.648 1.121 1.781 1.154 ;
      RECT 1.145 1.045 1.686 1.135 ;
      RECT 1.145 0.745 1.235 1.135 ;
      RECT 2.062 0.845 2.985 0.935 ;
      RECT 2.895 0.695 2.985 0.935 ;
      RECT 2.627 0.445 2.717 0.935 ;
      RECT 1.065 0.745 1.235 0.835 ;
      RECT 2.035 0.445 2.717 0.535 ;
      RECT 1.799 0.37 1.889 1.03 ;
      RECT 1.35 0.865 1.889 0.955 ;
      RECT 1.35 0.625 1.44 0.955 ;
      RECT 1.799 0.665 2.537 0.755 ;
      RECT 1.774 0.37 1.914 0.46 ;
      RECT 0.85 0.37 0.94 1.03 ;
      RECT 1.61 0.532 1.7 0.7 ;
      RECT 1.576 0.447 1.61 0.575 ;
      RECT 1.538 0.487 1.656 0.539 ;
      RECT 0.85 0.43 1.576 0.52 ;
      RECT 0.85 0.37 1.03 0.52 ;
  END
END DFFNX1H7R

MACRO DFFNX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNX2H7R 0 0 ;
  SIZE 5.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.4 1.48 ;
        RECT 5.087 0.92 5.227 1.48 ;
        RECT 4.572 1.225 4.712 1.48 ;
        RECT 3.732 1.225 3.872 1.48 ;
        RECT 2.289 1.095 2.429 1.48 ;
        RECT 1.47 1.225 1.61 1.48 ;
        RECT 0.31 1.12 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.4 0.08 ;
        RECT 4.522 -0.08 4.662 0.32 ;
        RECT 3.682 -0.08 3.822 0.34 ;
        RECT 2.305 -0.08 2.445 0.175 ;
        RECT 1.455 -0.08 1.595 0.16 ;
        RECT 0.36 -0.08 0.5 0.185 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.625 0.37 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.51 0.455 0.6 0.67 ;
        RECT 0.425 0.455 0.6 0.545 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.837 0.872 4.982 0.962 ;
        RECT 4.892 0.255 4.982 0.962 ;
        RECT 4.825 0.255 4.982 0.345 ;
      LAYER MET2 ;
        RECT 4.85 0.18 4.95 0.56 ;
      LAYER VIA1 ;
        RECT 4.855 0.255 4.945 0.345 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.077 0.865 4.217 1.04 ;
        RECT 3.715 0.865 4.217 0.955 ;
        RECT 3.715 0.455 4.062 0.545 ;
        RECT 3.972 0.33 4.062 0.545 ;
        RECT 3.715 0.455 3.805 0.955 ;
      LAYER MET2 ;
        RECT 3.85 0.23 3.95 0.76 ;
      LAYER VIA1 ;
        RECT 3.855 0.455 3.945 0.545 ;
    END
  END QN
  OBS
    LAYER MET1 ;
      RECT 4.005 1.14 4.436 1.23 ;
      RECT 3.994 1.096 4.005 1.225 ;
      RECT 3.994 1.14 4.482 1.207 ;
      RECT 3.948 1.068 3.994 1.196 ;
      RECT 4.398 1.121 4.512 1.169 ;
      RECT 3.91 1.121 4.043 1.154 ;
      RECT 3.092 1.045 3.948 1.135 ;
      RECT 4.436 1.079 4.558 1.131 ;
      RECT 4.482 1.041 4.512 1.169 ;
      RECT 4.512 0.587 4.602 1.086 ;
      RECT 3.092 0.404 3.182 1.135 ;
      RECT 4.512 0.587 4.802 0.727 ;
      RECT 2.809 0.404 3.182 0.494 ;
      RECT 4.332 0.32 4.422 0.987 ;
      RECT 3.897 0.645 4.422 0.735 ;
      RECT 4.207 0.32 4.422 0.41 ;
      RECT 0.585 1.14 1.055 1.23 ;
      RECT 0.585 0.94 0.675 1.23 ;
      RECT 0.07 0.94 0.675 1.03 ;
      RECT 0.07 0.275 0.16 1.03 ;
      RECT 3.362 0.17 3.452 0.816 ;
      RECT 0.07 0.275 0.681 0.365 ;
      RECT 0.591 0.17 0.681 0.365 ;
      RECT 2.229 0.265 2.609 0.355 ;
      RECT 2.218 0.221 2.229 0.35 ;
      RECT 1.377 0.25 1.671 0.34 ;
      RECT 2.218 0.265 2.655 0.332 ;
      RECT 2.172 0.193 2.218 0.321 ;
      RECT 1.335 0.25 1.713 0.319 ;
      RECT 1.297 0.25 1.751 0.279 ;
      RECT 2.571 0.246 2.704 0.279 ;
      RECT 2.655 0.175 2.666 0.304 ;
      RECT 2.134 0.246 2.267 0.279 ;
      RECT 2.666 0.17 3.452 0.26 ;
      RECT 1.713 0.17 2.172 0.26 ;
      RECT 1.671 0.191 1.713 0.319 ;
      RECT 0.591 0.231 1.415 0.26 ;
      RECT 2.609 0.204 3.452 0.26 ;
      RECT 1.633 0.231 2.229 0.26 ;
      RECT 0.591 0.191 1.377 0.26 ;
      RECT 0.591 0.17 1.335 0.26 ;
      RECT 1.743 1.14 2.152 1.23 ;
      RECT 2.062 0.845 2.152 1.23 ;
      RECT 1.732 1.096 1.743 1.225 ;
      RECT 1.686 1.068 1.732 1.196 ;
      RECT 1.648 1.121 1.781 1.154 ;
      RECT 1.145 1.045 1.686 1.135 ;
      RECT 1.145 0.745 1.235 1.135 ;
      RECT 2.062 0.845 2.985 0.935 ;
      RECT 2.895 0.655 2.985 0.935 ;
      RECT 2.629 0.445 2.719 0.935 ;
      RECT 1.065 0.745 1.235 0.835 ;
      RECT 2.035 0.445 2.719 0.535 ;
      RECT 2.035 0.429 2.175 0.535 ;
      RECT 1.799 0.37 1.889 1.03 ;
      RECT 1.35 0.865 1.889 0.955 ;
      RECT 1.35 0.625 1.44 0.955 ;
      RECT 1.799 0.665 2.539 0.755 ;
      RECT 1.774 0.37 1.914 0.46 ;
      RECT 0.85 0.37 0.94 1.03 ;
      RECT 1.61 0.532 1.7 0.7 ;
      RECT 1.576 0.447 1.61 0.575 ;
      RECT 1.538 0.487 1.656 0.539 ;
      RECT 0.85 0.43 1.576 0.52 ;
      RECT 0.85 0.37 1.03 0.52 ;
  END
END DFFNX2H7R

MACRO DFFNX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNX3H7R 0 0 ;
  SIZE 5.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.6 1.48 ;
        RECT 5.42 0.995 5.51 1.48 ;
        RECT 4.88 1.225 5.02 1.48 ;
        RECT 4.323 1.225 4.463 1.48 ;
        RECT 3.755 1.225 3.895 1.48 ;
        RECT 2.384 1.07 2.474 1.48 ;
        RECT 1.54 1.225 1.68 1.48 ;
        RECT 0.31 1.12 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.6 0.08 ;
        RECT 5.28 -0.08 5.37 0.365 ;
        RECT 4.775 -0.08 4.865 0.35 ;
        RECT 4.295 -0.08 4.385 0.415 ;
        RECT 3.755 -0.08 3.895 0.365 ;
        RECT 2.414 -0.08 2.504 0.2 ;
        RECT 1.525 -0.08 1.665 0.16 ;
        RECT 0.36 -0.08 0.5 0.185 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.625 0.37 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.51 0.455 0.6 0.67 ;
        RECT 0.425 0.455 0.6 0.545 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.145 0.872 5.29 0.962 ;
        RECT 5.2 0.455 5.29 0.962 ;
        RECT 5.025 0.455 5.29 0.545 ;
        RECT 5.025 0.3 5.115 0.545 ;
      LAYER MET2 ;
        RECT 5.05 0.23 5.15 0.76 ;
      LAYER VIA1 ;
        RECT 5.055 0.455 5.145 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.064 0.865 4.154 1.01 ;
        RECT 3.785 0.455 4.135 0.545 ;
        RECT 4.045 0.33 4.135 0.545 ;
        RECT 3.785 0.865 4.154 0.955 ;
        RECT 3.785 0.455 3.875 0.955 ;
      LAYER MET2 ;
        RECT 3.85 0.23 3.95 0.76 ;
      LAYER VIA1 ;
        RECT 3.855 0.455 3.945 0.545 ;
    END
  END QN
  OBS
    LAYER MET1 ;
      RECT 3.988 1.1 4.23 1.19 ;
      RECT 3.971 1.1 4.247 1.182 ;
      RECT 4.554 1.077 4.808 1.167 ;
      RECT 3.933 1.1 4.285 1.154 ;
      RECT 4.522 1.077 4.82 1.151 ;
      RECT 4.247 1.045 4.56 1.135 ;
      RECT 4.192 1.081 4.866 1.132 ;
      RECT 4.23 1.053 4.247 1.182 ;
      RECT 3.162 1.081 4.026 1.135 ;
      RECT 4.82 0.642 4.91 1.087 ;
      RECT 3.162 1.053 3.988 1.135 ;
      RECT 4.77 1.058 4.91 1.087 ;
      RECT 4.808 1.033 4.82 1.161 ;
      RECT 4.23 1.061 4.592 1.135 ;
      RECT 3.162 1.045 3.971 1.135 ;
      RECT 3.162 0.375 3.252 1.135 ;
      RECT 4.82 0.642 5.11 0.782 ;
      RECT 2.879 0.375 3.252 0.465 ;
      RECT 4.64 0.645 4.73 0.987 ;
      RECT 3.967 0.645 4.73 0.735 ;
      RECT 4.525 0.315 4.615 0.735 ;
      RECT 0.585 1.14 1.125 1.23 ;
      RECT 0.585 0.94 0.675 1.23 ;
      RECT 0.07 0.94 0.675 1.03 ;
      RECT 0.07 0.275 0.16 1.03 ;
      RECT 3.435 0.17 3.525 0.917 ;
      RECT 2.338 0.29 2.664 0.38 ;
      RECT 0.07 0.275 0.681 0.365 ;
      RECT 0.591 0.17 0.681 0.365 ;
      RECT 2.302 0.234 2.338 0.362 ;
      RECT 2.302 0.29 2.71 0.357 ;
      RECT 1.447 0.25 1.741 0.34 ;
      RECT 2.256 0.193 2.302 0.321 ;
      RECT 1.405 0.25 1.783 0.319 ;
      RECT 2.626 0.271 2.746 0.316 ;
      RECT 2.256 0.271 2.376 0.321 ;
      RECT 2.218 0.17 2.256 0.279 ;
      RECT 1.367 0.25 1.821 0.279 ;
      RECT 2.664 0.229 2.784 0.279 ;
      RECT 2.71 0.188 2.746 0.316 ;
      RECT 2.746 0.17 3.525 0.26 ;
      RECT 1.783 0.17 2.256 0.26 ;
      RECT 1.741 0.191 1.783 0.319 ;
      RECT 0.591 0.231 1.485 0.26 ;
      RECT 1.703 0.231 2.302 0.26 ;
      RECT 0.591 0.191 1.447 0.26 ;
      RECT 0.591 0.17 1.405 0.26 ;
      RECT 1.813 1.14 2.222 1.23 ;
      RECT 2.132 0.845 2.222 1.23 ;
      RECT 1.802 1.096 1.813 1.225 ;
      RECT 1.756 1.068 1.802 1.196 ;
      RECT 1.718 1.121 1.851 1.154 ;
      RECT 1.215 1.045 1.756 1.135 ;
      RECT 1.215 0.745 1.305 1.135 ;
      RECT 2.132 0.845 3.06 0.935 ;
      RECT 2.97 0.635 3.06 0.935 ;
      RECT 2.699 0.47 2.789 0.935 ;
      RECT 1.135 0.745 1.305 0.835 ;
      RECT 2.13 0.47 2.789 0.56 ;
      RECT 2.13 0.39 2.22 0.56 ;
      RECT 1.869 0.37 1.959 1.03 ;
      RECT 1.42 0.865 1.959 0.955 ;
      RECT 1.42 0.625 1.51 0.955 ;
      RECT 1.869 0.665 2.609 0.755 ;
      RECT 1.844 0.37 1.984 0.46 ;
      RECT 0.89 0.35 0.98 1.03 ;
      RECT 1.68 0.532 1.77 0.7 ;
      RECT 1.646 0.447 1.68 0.575 ;
      RECT 1.608 0.487 1.726 0.539 ;
      RECT 0.89 0.43 1.646 0.52 ;
      RECT 0.89 0.35 1.03 0.52 ;
  END
END DFFNX3H7R

MACRO DFFQX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFQX0P5H7R 0 0 ;
  SIZE 4.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.4 1.48 ;
        RECT 3.975 1.05 4.065 1.48 ;
        RECT 3.495 1.055 3.585 1.48 ;
        RECT 2.345 1.095 2.485 1.48 ;
        RECT 1.42 1.225 1.56 1.48 ;
        RECT 0.31 1.135 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.4 0.08 ;
        RECT 3.935 -0.08 4.075 0.21 ;
        RECT 3.305 -0.08 3.395 0.345 ;
        RECT 2.27 -0.08 2.41 0.16 ;
        RECT 1.43 -0.08 1.57 0.16 ;
        RECT 0.31 -0.08 0.45 0.325 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.585 0.35 0.855 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.425 0.575 0.65 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.225 0.275 4.345 1.045 ;
      LAYER MET2 ;
        RECT 4.25 0.625 4.35 1.16 ;
      LAYER VIA1 ;
        RECT 4.255 0.855 4.345 0.945 ;
    END
  END Q
  OBS
    LAYER MET1 ;
      RECT 3.7 0.93 3.874 1.02 ;
      RECT 3.7 0.93 3.92 0.997 ;
      RECT 3.836 0.911 3.966 0.951 ;
      RECT 3.874 0.869 3.966 0.951 ;
      RECT 3.874 0.869 4.012 0.905 ;
      RECT 3.92 0.823 4.02 0.878 ;
      RECT 3.966 0.777 4.066 0.851 ;
      RECT 4.012 0.75 4.02 0.878 ;
      RECT 4.02 0.3 4.11 0.806 ;
      RECT 3.485 0.3 3.575 0.525 ;
      RECT 3.485 0.3 4.11 0.39 ;
      RECT 2.96 1.095 3.405 1.185 ;
      RECT 3.315 0.615 3.405 1.185 ;
      RECT 3.315 0.615 3.93 0.705 ;
      RECT 3.297 0.576 3.315 0.704 ;
      RECT 3.251 0.544 3.297 0.672 ;
      RECT 3.205 0.498 3.251 0.626 ;
      RECT 3.205 0.6 3.345 0.626 ;
      RECT 3.159 0.452 3.205 0.58 ;
      RECT 3.113 0.406 3.159 0.534 ;
      RECT 3.067 0.36 3.113 0.488 ;
      RECT 3.021 0.314 3.067 0.442 ;
      RECT 2.975 0.268 3.021 0.396 ;
      RECT 2.937 0.314 3.067 0.354 ;
      RECT 2.82 0.245 2.975 0.335 ;
      RECT 2.054 1.067 2.144 1.23 ;
      RECT 2.1 1.022 2.19 1.105 ;
      RECT 2.144 0.977 2.267 1.024 ;
      RECT 2.19 0.934 2.229 1.063 ;
      RECT 3.135 0.762 3.225 1.005 ;
      RECT 2.229 0.915 3.225 1.005 ;
      RECT 3.12 0.686 3.135 0.815 ;
      RECT 3.074 0.656 3.12 0.784 ;
      RECT 3.074 0.717 3.181 0.784 ;
      RECT 3.028 0.61 3.074 0.738 ;
      RECT 2.982 0.564 3.028 0.692 ;
      RECT 2.936 0.518 2.982 0.646 ;
      RECT 2.898 0.564 3.028 0.604 ;
      RECT 2.635 0.495 2.936 0.585 ;
      RECT 2.635 0.281 2.725 0.585 ;
      RECT 2.015 0.281 2.725 0.371 ;
      RECT 1.352 0.25 1.646 0.34 ;
      RECT 1.31 0.25 1.688 0.319 ;
      RECT 2.015 0.17 2.105 0.371 ;
      RECT 1.272 0.25 1.726 0.279 ;
      RECT 1.688 0.17 2.105 0.26 ;
      RECT 1.608 0.231 2.105 0.26 ;
      RECT 1.646 0.191 1.688 0.319 ;
      RECT 1.04 0.231 1.39 0.26 ;
      RECT 1.04 0.191 1.352 0.26 ;
      RECT 1.04 0.17 1.31 0.26 ;
      RECT 0.71 1.12 1.16 1.21 ;
      RECT 1.07 1.015 1.16 1.21 ;
      RECT 0.71 0.485 0.8 1.21 ;
      RECT 1.07 1.015 1.911 1.105 ;
      RECT 1.07 1.015 1.957 1.082 ;
      RECT 0.07 0.955 0.8 1.045 ;
      RECT 1.873 0.996 2.003 1.036 ;
      RECT 1.911 0.954 2.003 1.036 ;
      RECT 0.07 0.275 0.16 1.045 ;
      RECT 1.957 0.908 2.049 0.99 ;
      RECT 2.003 0.862 2.095 0.944 ;
      RECT 2.003 0.862 2.141 0.898 ;
      RECT 2.049 0.816 2.163 0.864 ;
      RECT 2.095 0.77 2.201 0.834 ;
      RECT 2.141 0.736 2.163 0.864 ;
      RECT 2.163 0.725 2.849 0.815 ;
      RECT 1.305 0.835 1.835 0.925 ;
      RECT 1.78 0.37 1.87 0.908 ;
      RECT 1.305 0.745 1.445 0.925 ;
      RECT 1.78 0.515 2.545 0.605 ;
      RECT 1.78 0.37 1.885 0.605 ;
      RECT 1.745 0.37 1.885 0.46 ;
      RECT 0.89 0.365 0.98 1.03 ;
      RECT 1.383 0.54 1.69 0.63 ;
      RECT 1.338 0.479 1.383 0.608 ;
      RECT 1.292 0.434 1.338 0.562 ;
      RECT 1.292 0.521 1.421 0.562 ;
      RECT 1.246 0.388 1.292 0.516 ;
      RECT 1.208 0.434 1.338 0.474 ;
      RECT 0.89 0.365 1.246 0.455 ;
  END
END DFFQX0P5H7R

MACRO DFFQX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFQX1H7R 0 0 ;
  SIZE 4.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.4 1.48 ;
        RECT 3.96 1.06 4.1 1.48 ;
        RECT 3.49 1.055 3.58 1.48 ;
        RECT 2.345 1.095 2.485 1.48 ;
        RECT 1.42 1.225 1.56 1.48 ;
        RECT 0.31 1.135 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.4 0.08 ;
        RECT 3.985 -0.08 4.075 0.33 ;
        RECT 3.3 -0.08 3.39 0.33 ;
        RECT 2.245 -0.08 2.385 0.225 ;
        RECT 1.42 -0.08 1.56 0.16 ;
        RECT 0.31 -0.08 0.45 0.325 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.57 0.35 0.84 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.425 0.575 0.65 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.235 0.229 4.345 0.985 ;
      LAYER MET2 ;
        RECT 4.25 0.625 4.35 1.16 ;
      LAYER VIA1 ;
        RECT 4.255 0.855 4.345 0.945 ;
    END
  END Q
  OBS
    LAYER MET1 ;
      RECT 3.695 0.87 4.035 0.96 ;
      RECT 3.945 0.489 4.035 0.96 ;
      RECT 3.942 0.419 3.945 0.548 ;
      RECT 3.48 0.28 3.57 0.53 ;
      RECT 3.896 0.395 3.942 0.523 ;
      RECT 3.896 0.444 3.991 0.523 ;
      RECT 3.85 0.349 3.896 0.477 ;
      RECT 3.804 0.303 3.85 0.431 ;
      RECT 3.766 0.349 3.896 0.389 ;
      RECT 3.48 0.28 3.804 0.37 ;
      RECT 2.955 1.095 3.4 1.185 ;
      RECT 3.31 0.563 3.4 1.185 ;
      RECT 3.31 0.64 3.855 0.73 ;
      RECT 3.29 0.485 3.31 0.613 ;
      RECT 3.244 0.452 3.29 0.58 ;
      RECT 3.244 0.518 3.356 0.58 ;
      RECT 3.198 0.406 3.244 0.534 ;
      RECT 3.152 0.36 3.198 0.488 ;
      RECT 3.106 0.314 3.152 0.442 ;
      RECT 3.06 0.268 3.106 0.396 ;
      RECT 3.022 0.314 3.152 0.354 ;
      RECT 2.815 0.245 3.06 0.335 ;
      RECT 2.12 0.915 2.21 1.065 ;
      RECT 2.12 0.915 3.22 1.005 ;
      RECT 3.13 0.662 3.22 1.005 ;
      RECT 3.123 0.59 3.13 0.719 ;
      RECT 3.077 0.564 3.123 0.692 ;
      RECT 3.077 0.617 3.176 0.692 ;
      RECT 3.031 0.518 3.077 0.646 ;
      RECT 2.993 0.495 3.031 0.604 ;
      RECT 2.635 0.495 3.031 0.585 ;
      RECT 2.635 0.315 2.725 0.585 ;
      RECT 2.005 0.315 2.725 0.405 ;
      RECT 1.342 0.25 1.636 0.34 ;
      RECT 1.3 0.191 1.342 0.319 ;
      RECT 2.005 0.19 2.095 0.405 ;
      RECT 1.3 0.25 1.696 0.299 ;
      RECT 1.658 0.19 2.095 0.28 ;
      RECT 1.262 0.25 2.095 0.279 ;
      RECT 1.03 0.17 1.3 0.26 ;
      RECT 1.598 0.231 2.095 0.28 ;
      RECT 1.636 0.201 1.658 0.329 ;
      RECT 1.03 0.231 1.38 0.26 ;
      RECT 0.71 1.12 1.165 1.21 ;
      RECT 1.94 0.725 2.03 1.135 ;
      RECT 1.075 1.045 2.03 1.135 ;
      RECT 0.71 0.485 0.8 1.21 ;
      RECT 0.07 0.955 0.8 1.045 ;
      RECT 0.07 0.275 0.16 1.045 ;
      RECT 1.94 0.725 2.849 0.815 ;
      RECT 1.275 0.85 1.85 0.94 ;
      RECT 1.76 0.37 1.85 0.94 ;
      RECT 1.275 0.72 1.415 0.94 ;
      RECT 1.76 0.495 2.545 0.585 ;
      RECT 1.76 0.37 1.875 0.585 ;
      RECT 1.735 0.37 1.875 0.46 ;
      RECT 0.89 0.37 0.98 1.03 ;
      RECT 1.373 0.54 1.67 0.63 ;
      RECT 1.333 0.482 1.373 0.61 ;
      RECT 1.287 0.439 1.333 0.567 ;
      RECT 1.287 0.521 1.411 0.567 ;
      RECT 1.241 0.393 1.287 0.521 ;
      RECT 1.203 0.439 1.333 0.479 ;
      RECT 0.89 0.37 1.241 0.46 ;
  END
END DFFQX1H7R

MACRO DFFQX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFQX2H7R 0 0 ;
  SIZE 4.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.6 1.48 ;
        RECT 4.065 1.08 4.205 1.48 ;
        RECT 3.595 1.055 3.685 1.48 ;
        RECT 2.34 1.095 2.48 1.48 ;
        RECT 1.415 1.225 1.555 1.48 ;
        RECT 0.31 1.15 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.6 0.08 ;
        RECT 3.915 -0.08 4.055 0.21 ;
        RECT 3.37 -0.08 3.46 0.33 ;
        RECT 2.24 -0.08 2.38 0.215 ;
        RECT 1.4 -0.08 1.54 0.16 ;
        RECT 0.295 -0.08 0.435 0.325 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.565 0.35 0.835 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.42 0.575 0.645 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.34 0.255 4.43 1.145 ;
        RECT 4.225 0.255 4.43 0.345 ;
      LAYER MET2 ;
        RECT 4.25 0.18 4.35 0.56 ;
      LAYER VIA1 ;
        RECT 4.255 0.255 4.345 0.345 ;
    END
  END Q
  OBS
    LAYER MET1 ;
      RECT 3.8 0.895 4.125 0.985 ;
      RECT 4.035 0.3 4.125 0.985 ;
      RECT 3.595 0.3 3.685 0.625 ;
      RECT 3.595 0.3 4.125 0.39 ;
      RECT 2.954 1.095 3.505 1.185 ;
      RECT 3.415 0.575 3.505 1.185 ;
      RECT 3.415 0.715 3.945 0.805 ;
      RECT 3.855 0.625 3.945 0.805 ;
      RECT 3.383 0.491 3.415 0.619 ;
      RECT 3.337 0.452 3.383 0.58 ;
      RECT 3.337 0.53 3.461 0.58 ;
      RECT 3.291 0.406 3.337 0.534 ;
      RECT 3.245 0.36 3.291 0.488 ;
      RECT 3.199 0.314 3.245 0.442 ;
      RECT 3.153 0.268 3.199 0.396 ;
      RECT 3.115 0.314 3.245 0.354 ;
      RECT 2.825 0.245 3.153 0.335 ;
      RECT 2.115 0.915 2.205 1.055 ;
      RECT 2.115 0.915 3.325 1.005 ;
      RECT 3.235 0.661 3.325 1.005 ;
      RECT 3.193 0.572 3.235 0.7 ;
      RECT 3.193 0.616 3.281 0.7 ;
      RECT 3.147 0.528 3.193 0.656 ;
      RECT 3.109 0.572 3.235 0.614 ;
      RECT 2.645 0.505 3.147 0.595 ;
      RECT 2.645 0.306 2.735 0.595 ;
      RECT 1.985 0.306 2.735 0.396 ;
      RECT 1.307 0.25 1.616 0.34 ;
      RECT 1.265 0.25 1.658 0.319 ;
      RECT 1.985 0.17 2.075 0.396 ;
      RECT 1.227 0.25 1.696 0.279 ;
      RECT 1.658 0.17 2.075 0.26 ;
      RECT 1.578 0.231 2.075 0.26 ;
      RECT 1.616 0.191 1.658 0.319 ;
      RECT 1.01 0.231 1.345 0.26 ;
      RECT 1.01 0.191 1.307 0.26 ;
      RECT 1.01 0.17 1.265 0.26 ;
      RECT 0.705 1.12 1.155 1.21 ;
      RECT 1.935 0.705 2.025 1.135 ;
      RECT 1.065 1.045 2.025 1.135 ;
      RECT 0.705 0.485 0.795 1.21 ;
      RECT 0.07 0.955 0.795 1.045 ;
      RECT 0.07 0.275 0.16 1.045 ;
      RECT 1.935 0.705 3.09 0.795 ;
      RECT 1.27 0.85 1.845 0.94 ;
      RECT 1.755 0.37 1.845 0.94 ;
      RECT 1.27 0.72 1.41 0.94 ;
      RECT 1.755 0.515 2.546 0.605 ;
      RECT 1.755 0.37 1.855 0.605 ;
      RECT 1.715 0.37 1.855 0.46 ;
      RECT 0.885 0.37 0.975 1.03 ;
      RECT 1.338 0.54 1.665 0.63 ;
      RECT 1.298 0.482 1.338 0.61 ;
      RECT 1.252 0.439 1.298 0.567 ;
      RECT 1.252 0.521 1.376 0.567 ;
      RECT 1.206 0.393 1.252 0.521 ;
      RECT 1.168 0.439 1.298 0.479 ;
      RECT 0.885 0.37 1.206 0.46 ;
  END
END DFFQX2H7R

MACRO DFFQX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFQX3H7R 0 0 ;
  SIZE 4.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.8 1.48 ;
        RECT 4.595 1.035 4.685 1.48 ;
        RECT 4.095 1.05 4.185 1.48 ;
        RECT 3.6 1.055 3.69 1.48 ;
        RECT 2.405 1.095 2.545 1.48 ;
        RECT 1.48 1.225 1.62 1.48 ;
        RECT 0.31 1.105 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.8 0.08 ;
        RECT 4.525 -0.08 4.615 0.355 ;
        RECT 3.92 -0.08 4.06 0.21 ;
        RECT 3.373 -0.08 3.463 0.33 ;
        RECT 2.305 -0.08 2.445 0.215 ;
        RECT 1.465 -0.08 1.605 0.16 ;
        RECT 0.295 -0.08 0.435 0.325 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.535 0.35 0.805 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.42 0.575 0.645 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.345 0.255 4.435 1.01 ;
        RECT 4.225 0.255 4.435 0.345 ;
      LAYER MET2 ;
        RECT 4.25 0.18 4.35 0.56 ;
      LAYER VIA1 ;
        RECT 4.255 0.255 4.345 0.345 ;
    END
  END Q
  OBS
    LAYER MET1 ;
      RECT 3.805 0.93 3.994 1.02 ;
      RECT 4.04 0.3 4.086 0.951 ;
      RECT 3.956 0.911 4.086 0.951 ;
      RECT 3.994 0.869 4.04 0.997 ;
      RECT 4.04 0.3 4.13 0.906 ;
      RECT 3.6 0.3 3.69 0.625 ;
      RECT 3.6 0.3 4.13 0.39 ;
      RECT 3.065 1.095 3.51 1.185 ;
      RECT 3.42 0.573 3.51 1.185 ;
      RECT 3.42 0.715 3.95 0.805 ;
      RECT 3.86 0.625 3.95 0.805 ;
      RECT 3.39 0.49 3.42 0.618 ;
      RECT 3.344 0.452 3.39 0.58 ;
      RECT 3.344 0.528 3.466 0.58 ;
      RECT 3.298 0.406 3.344 0.534 ;
      RECT 3.252 0.36 3.298 0.488 ;
      RECT 3.206 0.314 3.252 0.442 ;
      RECT 3.16 0.268 3.206 0.396 ;
      RECT 3.122 0.314 3.252 0.354 ;
      RECT 2.885 0.245 3.16 0.335 ;
      RECT 2.18 0.915 2.27 1.08 ;
      RECT 2.18 0.915 3.33 1.005 ;
      RECT 3.24 0.666 3.33 1.005 ;
      RECT 3.239 0.597 3.24 0.726 ;
      RECT 3.193 0.574 3.239 0.702 ;
      RECT 3.193 0.621 3.286 0.702 ;
      RECT 3.147 0.528 3.193 0.656 ;
      RECT 3.109 0.505 3.147 0.614 ;
      RECT 2.705 0.505 3.147 0.595 ;
      RECT 2.705 0.305 2.795 0.595 ;
      RECT 2.05 0.305 2.795 0.395 ;
      RECT 1.387 0.25 1.681 0.34 ;
      RECT 1.345 0.191 1.387 0.319 ;
      RECT 2.05 0.19 2.14 0.395 ;
      RECT 1.345 0.25 1.741 0.299 ;
      RECT 1.703 0.19 2.14 0.28 ;
      RECT 1.307 0.25 2.14 0.279 ;
      RECT 1.045 0.17 1.345 0.26 ;
      RECT 1.643 0.231 2.14 0.28 ;
      RECT 1.681 0.201 1.703 0.329 ;
      RECT 1.045 0.231 1.425 0.26 ;
      RECT 0.74 1.115 1.215 1.205 ;
      RECT 2 0.735 2.09 1.135 ;
      RECT 1.125 1.045 2.09 1.135 ;
      RECT 0.74 0.515 0.83 1.205 ;
      RECT 0.07 0.925 0.83 1.015 ;
      RECT 0.07 0.295 0.16 1.015 ;
      RECT 2 0.735 3.095 0.825 ;
      RECT 1.335 0.85 1.91 0.94 ;
      RECT 1.82 0.37 1.91 0.94 ;
      RECT 1.335 0.72 1.475 0.94 ;
      RECT 1.82 0.485 2.615 0.575 ;
      RECT 1.82 0.37 1.92 0.575 ;
      RECT 1.78 0.37 1.92 0.46 ;
      RECT 0.92 0.365 1.01 1 ;
      RECT 1.418 0.54 1.73 0.63 ;
      RECT 1.373 0.479 1.418 0.608 ;
      RECT 1.327 0.434 1.373 0.562 ;
      RECT 1.327 0.521 1.456 0.562 ;
      RECT 1.281 0.388 1.327 0.516 ;
      RECT 1.243 0.434 1.373 0.474 ;
      RECT 0.92 0.365 1.281 0.455 ;
  END
END DFFQX3H7R

MACRO DFFRQNX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRQNX1H7R 0 0 ;
  SIZE 5.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.6 1.48 ;
        RECT 5.378 1.055 5.468 1.48 ;
        RECT 4.608 1.225 4.748 1.48 ;
        RECT 2.864 1.225 3.004 1.48 ;
        RECT 2.324 1.225 2.464 1.48 ;
        RECT 1.164 1.225 1.304 1.48 ;
        RECT 0.31 1.225 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.6 0.08 ;
        RECT 5.032 -0.08 5.122 0.35 ;
        RECT 3.131 -0.08 3.271 0.175 ;
        RECT 2.299 -0.08 2.389 0.2 ;
        RECT 1.164 -0.08 1.304 0.175 ;
        RECT 0.31 -0.08 0.45 0.325 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.595 0.345 0.853 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.815 0.684 1.032 0.775 ;
        RECT 0.815 0.607 0.955 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.128 0.85 5.545 0.94 ;
        RECT 5.44 0.425 5.545 0.94 ;
        RECT 5.282 0.425 5.545 0.53 ;
        RECT 5.282 0.224 5.372 0.53 ;
        RECT 5.128 0.85 5.218 1.1 ;
      LAYER MET2 ;
        RECT 5.45 0.225 5.55 0.76 ;
      LAYER VIA1 ;
        RECT 5.455 0.455 5.545 0.545 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.804 0.655 3.092 0.806 ;
      LAYER MET2 ;
        RECT 2.85 0.43 2.95 0.96 ;
      LAYER VIA1 ;
        RECT 2.855 0.655 2.945 0.745 ;
    END
  END RN
  OBS
    LAYER MET1 ;
      RECT 4.865 1.035 4.997 1.175 ;
      RECT 4.907 0.445 4.997 1.175 ;
      RECT 4.907 0.62 5.297 0.71 ;
      RECT 4.442 0.445 4.582 0.61 ;
      RECT 4.442 0.445 4.997 0.535 ;
      RECT 4.782 0.225 4.872 0.535 ;
      RECT 3.747 0.843 3.837 1.015 ;
      RECT 3.747 0.843 3.883 0.881 ;
      RECT 3.793 0.798 3.898 0.851 ;
      RECT 3.793 0.798 3.936 0.824 ;
      RECT 4.727 0.635 4.817 0.805 ;
      RECT 3.837 0.753 4.817 0.805 ;
      RECT 3.898 0.715 4.817 0.805 ;
      RECT 3.883 0.722 4.817 0.805 ;
      RECT 4.062 0.35 4.152 0.805 ;
      RECT 4.037 0.35 4.177 0.44 ;
      RECT 3.144 1.14 4.127 1.23 ;
      RECT 4.037 0.9 4.127 1.23 ;
      RECT 3.144 1.107 3.284 1.23 ;
      RECT 4.037 0.9 4.457 0.99 ;
      RECT 3.432 0.605 3.522 1.005 ;
      RECT 2.624 0.47 2.714 0.991 ;
      RECT 3.432 0.605 3.79 0.695 ;
      RECT 3.432 0.605 3.857 0.651 ;
      RECT 3.388 0.513 3.432 0.641 ;
      RECT 3.811 0.35 3.901 0.606 ;
      RECT 3.752 0.586 3.901 0.606 ;
      RECT 3.79 0.556 3.811 0.685 ;
      RECT 3.388 0.593 3.502 0.641 ;
      RECT 3.342 0.468 3.388 0.596 ;
      RECT 3.342 0.558 3.478 0.596 ;
      RECT 3.329 0.558 3.478 0.567 ;
      RECT 2.634 0.445 3.342 0.56 ;
      RECT 2.189 0.47 3.388 0.56 ;
      RECT 2.634 0.35 2.774 0.56 ;
      RECT 3.786 0.35 3.926 0.44 ;
      RECT 0.57 0.865 0.765 0.955 ;
      RECT 0.635 0.17 0.725 0.955 ;
      RECT 1.929 0.48 2.069 0.57 ;
      RECT 3.581 0.375 3.671 0.515 ;
      RECT 1.954 0.17 2.044 0.57 ;
      RECT 3.49 0.375 3.671 0.465 ;
      RECT 3.464 0.324 3.49 0.452 ;
      RECT 3.418 0.288 3.464 0.416 ;
      RECT 1.954 0.29 2.465 0.38 ;
      RECT 3.418 0.356 3.528 0.416 ;
      RECT 3.38 0.265 3.418 0.374 ;
      RECT 1.954 0.29 2.511 0.357 ;
      RECT 2.932 0.265 3.418 0.355 ;
      RECT 1.088 0.265 1.38 0.355 ;
      RECT 1.077 0.221 1.088 0.35 ;
      RECT 0.575 0.26 0.725 0.35 ;
      RECT 1.077 0.265 1.426 0.332 ;
      RECT 1.031 0.193 1.077 0.321 ;
      RECT 2.427 0.271 2.547 0.316 ;
      RECT 2.465 0.229 2.585 0.279 ;
      RECT 2.511 0.188 2.547 0.316 ;
      RECT 2.932 0.17 3.022 0.355 ;
      RECT 1.342 0.246 1.475 0.279 ;
      RECT 1.426 0.175 1.437 0.304 ;
      RECT 0.993 0.246 1.126 0.279 ;
      RECT 2.547 0.17 3.022 0.26 ;
      RECT 1.437 0.17 2.044 0.26 ;
      RECT 0.635 0.17 1.031 0.26 ;
      RECT 1.38 0.204 2.044 0.26 ;
      RECT 1.464 1.14 2.094 1.23 ;
      RECT 2.004 0.85 2.094 1.23 ;
      RECT 2.549 1.092 2.779 1.182 ;
      RECT 2.54 1.049 2.549 1.178 ;
      RECT 2.502 1.092 2.807 1.154 ;
      RECT 1.464 0.62 1.554 1.23 ;
      RECT 2.004 1.045 2.54 1.135 ;
      RECT 0.148 1.045 1.554 1.135 ;
      RECT 2.741 1.073 2.853 1.131 ;
      RECT 2.779 1.04 2.807 1.168 ;
      RECT 2.004 1.073 2.587 1.135 ;
      RECT 2.807 0.915 2.897 1.086 ;
      RECT 0.148 0.943 0.238 1.135 ;
      RECT 0.045 0.943 0.238 1.033 ;
      RECT 2.807 0.915 3.33 1.005 ;
      RECT 3.24 0.722 3.33 1.005 ;
      RECT 0.045 0.265 0.135 1.033 ;
      RECT 1.979 0.85 2.119 0.94 ;
      RECT 0.455 0.479 0.545 0.758 ;
      RECT 1.464 0.62 1.654 0.71 ;
      RECT 1.564 0.545 1.654 0.71 ;
      RECT 0.424 0.479 0.545 0.521 ;
      RECT 0.045 0.415 0.462 0.505 ;
      RECT 0.045 0.438 0.508 0.505 ;
      RECT 0.045 0.265 0.185 0.505 ;
      RECT 1.704 0.96 1.844 1.05 ;
      RECT 1.744 0.67 1.844 1.05 ;
      RECT 2.444 0.67 2.534 0.835 ;
      RECT 1.744 0.67 2.534 0.76 ;
      RECT 1.744 0.35 1.834 1.05 ;
      RECT 1.694 0.35 1.834 0.44 ;
      RECT 0.884 0.865 1.364 0.955 ;
      RECT 1.274 0.621 1.364 0.955 ;
      RECT 1.188 0.621 1.364 0.711 ;
      RECT 1.17 0.574 1.188 0.702 ;
      RECT 1.124 0.542 1.17 0.67 ;
      RECT 1.078 0.496 1.124 0.624 ;
      RECT 1.078 0.602 1.226 0.624 ;
      RECT 1.032 0.45 1.078 0.578 ;
      RECT 0.994 0.496 1.124 0.536 ;
      RECT 0.815 0.427 1.032 0.517 ;
      RECT 0.815 0.35 0.955 0.517 ;
      RECT 3.541 0.17 4.667 0.26 ;
  END
END DFFRQNX1H7R

MACRO DFFRQNX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRQNX2H7R 0 0 ;
  SIZE 5.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.8 1.48 ;
        RECT 5.415 1.225 5.555 1.48 ;
        RECT 4.608 1.225 4.748 1.48 ;
        RECT 2.864 1.225 3.004 1.48 ;
        RECT 2.324 1.225 2.464 1.48 ;
        RECT 1.164 1.225 1.304 1.48 ;
        RECT 0.31 1.225 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.8 0.08 ;
        RECT 5.532 -0.08 5.622 0.35 ;
        RECT 5.032 -0.08 5.122 0.35 ;
        RECT 3.131 -0.08 3.271 0.175 ;
        RECT 2.299 -0.08 2.389 0.2 ;
        RECT 1.164 -0.08 1.304 0.175 ;
        RECT 0.31 -0.08 0.45 0.325 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.595 0.345 0.853 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.815 0.684 1.032 0.775 ;
        RECT 0.815 0.607 0.955 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.1 0.85 5.575 0.94 ;
        RECT 5.425 0.44 5.575 0.94 ;
        RECT 5.282 0.44 5.575 0.53 ;
        RECT 5.282 0.224 5.372 0.53 ;
      LAYER MET2 ;
        RECT 5.45 0.225 5.55 0.76 ;
      LAYER VIA1 ;
        RECT 5.455 0.455 5.545 0.545 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.804 0.655 3.092 0.806 ;
      LAYER MET2 ;
        RECT 2.85 0.43 2.95 0.96 ;
      LAYER VIA1 ;
        RECT 2.855 0.655 2.945 0.745 ;
    END
  END RN
  OBS
    LAYER MET1 ;
      RECT 4.875 1.035 4.997 1.175 ;
      RECT 4.907 0.445 4.997 1.175 ;
      RECT 4.907 0.62 5.297 0.71 ;
      RECT 4.442 0.445 4.582 0.61 ;
      RECT 4.442 0.445 4.997 0.535 ;
      RECT 4.782 0.24 4.872 0.535 ;
      RECT 3.747 0.843 3.837 1.015 ;
      RECT 3.747 0.843 3.883 0.881 ;
      RECT 3.793 0.798 3.898 0.851 ;
      RECT 3.793 0.798 3.936 0.824 ;
      RECT 4.727 0.635 4.817 0.805 ;
      RECT 3.837 0.753 4.817 0.805 ;
      RECT 3.898 0.715 4.817 0.805 ;
      RECT 3.883 0.722 4.817 0.805 ;
      RECT 4.062 0.35 4.152 0.805 ;
      RECT 4.037 0.35 4.177 0.44 ;
      RECT 3.144 1.14 4.127 1.23 ;
      RECT 4.037 0.9 4.127 1.23 ;
      RECT 3.144 1.107 3.284 1.23 ;
      RECT 4.037 0.9 4.457 0.99 ;
      RECT 3.432 0.605 3.522 1.005 ;
      RECT 2.624 0.388 2.714 0.991 ;
      RECT 3.432 0.605 3.79 0.695 ;
      RECT 3.432 0.605 3.857 0.651 ;
      RECT 3.388 0.513 3.432 0.641 ;
      RECT 3.811 0.35 3.901 0.606 ;
      RECT 3.752 0.586 3.901 0.606 ;
      RECT 3.79 0.556 3.811 0.685 ;
      RECT 3.388 0.593 3.502 0.641 ;
      RECT 3.342 0.468 3.388 0.596 ;
      RECT 3.342 0.558 3.478 0.596 ;
      RECT 2.189 0.47 2.745 0.56 ;
      RECT 3.304 0.513 3.432 0.554 ;
      RECT 2.605 0.445 3.342 0.535 ;
      RECT 2.605 0.388 2.774 0.535 ;
      RECT 2.634 0.35 2.774 0.535 ;
      RECT 3.786 0.35 3.926 0.44 ;
      RECT 0.57 0.865 0.73 0.955 ;
      RECT 0.635 0.17 0.725 0.955 ;
      RECT 1.929 0.48 2.069 0.57 ;
      RECT 3.581 0.375 3.671 0.515 ;
      RECT 1.954 0.17 2.044 0.57 ;
      RECT 3.49 0.375 3.671 0.465 ;
      RECT 3.464 0.324 3.49 0.452 ;
      RECT 3.418 0.288 3.464 0.416 ;
      RECT 1.954 0.29 2.465 0.38 ;
      RECT 3.418 0.356 3.528 0.416 ;
      RECT 3.38 0.265 3.418 0.374 ;
      RECT 1.954 0.29 2.511 0.357 ;
      RECT 2.932 0.265 3.418 0.355 ;
      RECT 1.088 0.265 1.38 0.355 ;
      RECT 1.077 0.221 1.088 0.35 ;
      RECT 0.575 0.26 0.725 0.35 ;
      RECT 1.077 0.265 1.426 0.332 ;
      RECT 1.031 0.193 1.077 0.321 ;
      RECT 2.427 0.271 2.547 0.316 ;
      RECT 2.465 0.229 2.585 0.279 ;
      RECT 2.511 0.188 2.547 0.316 ;
      RECT 2.932 0.17 3.022 0.355 ;
      RECT 1.342 0.246 1.475 0.279 ;
      RECT 1.426 0.175 1.437 0.304 ;
      RECT 0.993 0.246 1.126 0.279 ;
      RECT 2.547 0.17 3.022 0.26 ;
      RECT 1.437 0.17 2.044 0.26 ;
      RECT 0.635 0.17 1.031 0.26 ;
      RECT 1.38 0.204 2.044 0.26 ;
      RECT 1.464 1.14 2.094 1.23 ;
      RECT 2.004 0.85 2.094 1.23 ;
      RECT 2.549 1.092 2.779 1.182 ;
      RECT 2.54 1.049 2.549 1.178 ;
      RECT 2.502 1.092 2.807 1.154 ;
      RECT 1.464 0.62 1.554 1.23 ;
      RECT 2.004 1.045 2.54 1.135 ;
      RECT 0.148 1.045 1.554 1.135 ;
      RECT 2.741 1.073 2.853 1.131 ;
      RECT 2.779 1.04 2.807 1.168 ;
      RECT 2.004 1.073 2.587 1.135 ;
      RECT 2.807 0.915 2.897 1.086 ;
      RECT 0.148 0.943 0.238 1.135 ;
      RECT 0.045 0.943 0.238 1.033 ;
      RECT 2.807 0.915 3.33 1.005 ;
      RECT 3.24 0.722 3.33 1.005 ;
      RECT 0.045 0.265 0.135 1.033 ;
      RECT 1.979 0.85 2.119 0.94 ;
      RECT 0.455 0.479 0.545 0.758 ;
      RECT 1.464 0.62 1.654 0.71 ;
      RECT 1.564 0.545 1.654 0.71 ;
      RECT 0.424 0.479 0.545 0.521 ;
      RECT 0.045 0.415 0.462 0.505 ;
      RECT 0.045 0.438 0.508 0.505 ;
      RECT 0.045 0.265 0.185 0.505 ;
      RECT 1.704 0.96 1.844 1.05 ;
      RECT 1.744 0.35 1.834 1.05 ;
      RECT 2.444 0.67 2.534 0.835 ;
      RECT 1.744 0.67 2.534 0.76 ;
      RECT 1.694 0.35 1.834 0.44 ;
      RECT 0.884 0.865 1.364 0.955 ;
      RECT 1.274 0.621 1.364 0.955 ;
      RECT 1.188 0.621 1.364 0.711 ;
      RECT 1.17 0.574 1.188 0.702 ;
      RECT 1.124 0.542 1.17 0.67 ;
      RECT 1.078 0.496 1.124 0.624 ;
      RECT 1.078 0.602 1.226 0.624 ;
      RECT 1.032 0.45 1.078 0.578 ;
      RECT 0.994 0.496 1.124 0.536 ;
      RECT 0.855 0.427 1.032 0.517 ;
      RECT 0.815 0.35 0.955 0.44 ;
      RECT 3.541 0.17 4.667 0.26 ;
  END
END DFFRQNX2H7R

MACRO DFFRQX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRQX0P5H7R 0 0 ;
  SIZE 5.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.6 1.48 ;
        RECT 5.128 1.005 5.218 1.48 ;
        RECT 4.608 1.225 4.748 1.48 ;
        RECT 2.864 1.225 3.004 1.48 ;
        RECT 2.324 1.225 2.464 1.48 ;
        RECT 1.164 1.225 1.304 1.48 ;
        RECT 0.31 1.225 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.6 0.08 ;
        RECT 5.128 -0.08 5.218 0.374 ;
        RECT 3.131 -0.08 3.271 0.175 ;
        RECT 2.299 -0.08 2.389 0.2 ;
        RECT 1.164 -0.08 1.304 0.175 ;
        RECT 0.335 -0.08 0.425 0.245 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.59 0.345 0.815 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.815 0.679 0.992 0.775 ;
        RECT 0.815 0.607 0.955 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.378 0.284 5.468 1.015 ;
        RECT 5.225 0.655 5.468 0.745 ;
      LAYER MET2 ;
        RECT 5.25 0.425 5.35 0.96 ;
      LAYER VIA1 ;
        RECT 5.255 0.655 5.345 0.745 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.995 0.625 3.145 0.805 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END RN
  OBS
    LAYER MET1 ;
      RECT 4.898 0.895 4.988 1.123 ;
      RECT 4.928 0.52 5.018 0.985 ;
      RECT 4.433 0.52 5.018 0.61 ;
      RECT 4.878 0.284 4.968 0.61 ;
      RECT 3.144 1.107 4.506 1.197 ;
      RECT 4.468 1.088 4.593 1.133 ;
      RECT 4.506 1.048 4.547 1.177 ;
      RECT 3.707 1.03 3.847 1.197 ;
      RECT 4.547 0.715 4.637 1.088 ;
      RECT 4.087 0.715 4.838 0.805 ;
      RECT 4.087 0.35 4.177 0.805 ;
      RECT 4.037 0.35 4.177 0.44 ;
      RECT 2.624 0.47 2.714 0.991 ;
      RECT 3.432 0.85 3.855 0.94 ;
      RECT 3.765 0.35 3.855 0.94 ;
      RECT 3.5 0.641 3.855 0.731 ;
      RECT 3.48 0.593 3.5 0.721 ;
      RECT 3.434 0.56 3.48 0.688 ;
      RECT 3.388 0.514 3.434 0.642 ;
      RECT 3.388 0.622 3.538 0.642 ;
      RECT 3.342 0.468 3.388 0.596 ;
      RECT 2.189 0.47 2.714 0.56 ;
      RECT 3.304 0.514 3.434 0.554 ;
      RECT 2.634 0.445 3.342 0.535 ;
      RECT 2.634 0.35 2.774 0.535 ;
      RECT 3.765 0.35 3.926 0.44 ;
      RECT 0.57 0.865 0.725 0.955 ;
      RECT 0.635 0.17 0.725 0.955 ;
      RECT 1.929 0.48 2.069 0.57 ;
      RECT 1.979 0.17 2.069 0.57 ;
      RECT 3.581 0.41 3.671 0.55 ;
      RECT 3.525 0.41 3.671 0.5 ;
      RECT 3.51 0.364 3.525 0.493 ;
      RECT 3.464 0.334 3.51 0.462 ;
      RECT 3.418 0.288 3.464 0.416 ;
      RECT 3.418 0.391 3.563 0.416 ;
      RECT 1.979 0.29 2.465 0.38 ;
      RECT 0.575 0.285 0.725 0.375 ;
      RECT 3.38 0.265 3.418 0.374 ;
      RECT 1.979 0.29 2.511 0.357 ;
      RECT 2.932 0.265 3.418 0.355 ;
      RECT 1.088 0.265 1.38 0.355 ;
      RECT 1.077 0.221 1.088 0.35 ;
      RECT 1.077 0.265 1.426 0.332 ;
      RECT 1.031 0.193 1.077 0.321 ;
      RECT 2.427 0.271 2.547 0.316 ;
      RECT 2.465 0.229 2.585 0.279 ;
      RECT 2.511 0.188 2.547 0.316 ;
      RECT 2.932 0.17 3.022 0.355 ;
      RECT 1.342 0.246 1.475 0.279 ;
      RECT 1.426 0.175 1.437 0.304 ;
      RECT 0.993 0.246 1.126 0.279 ;
      RECT 2.547 0.17 3.022 0.26 ;
      RECT 1.437 0.17 2.069 0.26 ;
      RECT 0.635 0.17 1.031 0.26 ;
      RECT 1.38 0.204 2.069 0.26 ;
      RECT 1.464 1.115 2.119 1.205 ;
      RECT 2.029 0.85 2.119 1.205 ;
      RECT 2.549 1.092 2.779 1.182 ;
      RECT 2.54 1.049 2.549 1.178 ;
      RECT 2.54 1.092 2.825 1.159 ;
      RECT 2.502 1.092 2.825 1.154 ;
      RECT 2.029 1.045 2.54 1.135 ;
      RECT 0.148 1.045 1.554 1.135 ;
      RECT 1.464 0.62 1.554 1.205 ;
      RECT 2.741 1.073 2.871 1.113 ;
      RECT 2.029 1.073 2.587 1.135 ;
      RECT 2.779 1.031 2.871 1.113 ;
      RECT 0.148 0.943 0.238 1.135 ;
      RECT 0.045 0.943 0.238 1.033 ;
      RECT 2.825 0.985 2.918 1.044 ;
      RECT 2.871 0.939 2.917 1.067 ;
      RECT 2.825 0.985 2.956 1.024 ;
      RECT 3.252 0.702 3.342 1.005 ;
      RECT 2.917 0.915 3.342 1.005 ;
      RECT 0.045 0.335 0.135 1.033 ;
      RECT 1.979 0.85 2.119 0.94 ;
      RECT 1.464 0.62 1.654 0.71 ;
      RECT 1.564 0.545 1.654 0.71 ;
      RECT 0.455 0.476 0.545 0.66 ;
      RECT 0.428 0.394 0.455 0.523 ;
      RECT 0.382 0.358 0.428 0.486 ;
      RECT 0.382 0.431 0.501 0.486 ;
      RECT 0.344 0.335 0.382 0.444 ;
      RECT 0.045 0.335 0.382 0.425 ;
      RECT 1.669 0.935 1.834 1.025 ;
      RECT 1.744 0.35 1.834 1.025 ;
      RECT 2.444 0.67 2.534 0.821 ;
      RECT 1.744 0.67 2.534 0.76 ;
      RECT 1.694 0.35 1.834 0.44 ;
      RECT 0.884 0.865 1.364 0.955 ;
      RECT 1.274 0.621 1.364 0.955 ;
      RECT 1.188 0.621 1.364 0.711 ;
      RECT 1.185 0.581 1.188 0.71 ;
      RECT 1.139 0.557 1.185 0.685 ;
      RECT 1.093 0.511 1.139 0.639 ;
      RECT 1.093 0.602 1.226 0.639 ;
      RECT 1.047 0.465 1.093 0.593 ;
      RECT 1.001 0.419 1.047 0.547 ;
      RECT 0.955 0.373 1.001 0.501 ;
      RECT 0.917 0.419 1.047 0.459 ;
      RECT 0.815 0.35 0.955 0.44 ;
      RECT 3.541 0.17 4.667 0.26 ;
      RECT 4.037 0.9 4.457 0.99 ;
  END
END DFFRQX0P5H7R

MACRO DFFRQX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRQX1H7R 0 0 ;
  SIZE 5.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.6 1.48 ;
        RECT 5.128 1.055 5.218 1.48 ;
        RECT 4.608 1.225 4.748 1.48 ;
        RECT 2.864 1.225 3.004 1.48 ;
        RECT 2.324 1.225 2.464 1.48 ;
        RECT 1.164 1.225 1.304 1.48 ;
        RECT 0.31 1.225 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.6 0.08 ;
        RECT 5.128 -0.08 5.218 0.354 ;
        RECT 3.131 -0.08 3.271 0.175 ;
        RECT 2.299 -0.08 2.389 0.2 ;
        RECT 1.164 -0.08 1.304 0.175 ;
        RECT 0.335 -0.08 0.425 0.245 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.585 0.345 0.81 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.815 0.639 0.982 0.775 ;
        RECT 0.815 0.607 0.955 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.378 0.284 5.468 1.015 ;
        RECT 5.225 0.655 5.468 0.745 ;
      LAYER MET2 ;
        RECT 5.25 0.425 5.35 0.96 ;
      LAYER VIA1 ;
        RECT 5.255 0.655 5.345 0.745 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.995 0.625 3.145 0.805 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END RN
  OBS
    LAYER MET1 ;
      RECT 4.873 0.9 5.018 0.99 ;
      RECT 4.928 0.52 5.018 0.99 ;
      RECT 4.442 0.52 5.018 0.61 ;
      RECT 4.878 0.284 4.968 0.61 ;
      RECT 3.144 1.14 4.473 1.23 ;
      RECT 3.144 1.14 4.519 1.207 ;
      RECT 4.435 1.121 4.547 1.17 ;
      RECT 3.707 1.03 3.847 1.23 ;
      RECT 3.144 1.107 3.284 1.23 ;
      RECT 4.473 1.079 4.593 1.133 ;
      RECT 4.519 1.042 4.547 1.17 ;
      RECT 4.547 0.715 4.637 1.088 ;
      RECT 4.087 0.715 4.838 0.805 ;
      RECT 4.087 0.35 4.177 0.805 ;
      RECT 4.037 0.35 4.177 0.44 ;
      RECT 2.624 0.47 2.714 0.991 ;
      RECT 3.432 0.85 3.876 0.94 ;
      RECT 3.786 0.35 3.876 0.94 ;
      RECT 3.5 0.641 3.876 0.731 ;
      RECT 3.48 0.593 3.5 0.721 ;
      RECT 3.434 0.56 3.48 0.688 ;
      RECT 3.388 0.514 3.434 0.642 ;
      RECT 3.388 0.622 3.538 0.642 ;
      RECT 3.342 0.468 3.388 0.596 ;
      RECT 2.189 0.47 2.714 0.56 ;
      RECT 3.304 0.514 3.434 0.554 ;
      RECT 2.634 0.445 3.342 0.535 ;
      RECT 2.634 0.35 2.774 0.535 ;
      RECT 3.786 0.35 3.926 0.44 ;
      RECT 0.57 0.865 0.725 0.955 ;
      RECT 0.635 0.17 0.725 0.955 ;
      RECT 1.929 0.48 2.069 0.57 ;
      RECT 3.581 0.375 3.671 0.515 ;
      RECT 1.954 0.17 2.044 0.57 ;
      RECT 3.49 0.375 3.671 0.465 ;
      RECT 3.464 0.324 3.49 0.452 ;
      RECT 3.418 0.288 3.464 0.416 ;
      RECT 1.954 0.29 2.465 0.38 ;
      RECT 0.575 0.285 0.725 0.375 ;
      RECT 3.418 0.356 3.528 0.416 ;
      RECT 3.38 0.265 3.418 0.374 ;
      RECT 1.954 0.29 2.511 0.357 ;
      RECT 2.932 0.265 3.418 0.355 ;
      RECT 1.088 0.265 1.38 0.355 ;
      RECT 1.077 0.221 1.088 0.35 ;
      RECT 1.077 0.265 1.426 0.332 ;
      RECT 1.031 0.193 1.077 0.321 ;
      RECT 2.427 0.271 2.547 0.316 ;
      RECT 2.465 0.229 2.585 0.279 ;
      RECT 2.511 0.188 2.547 0.316 ;
      RECT 2.932 0.17 3.022 0.355 ;
      RECT 1.342 0.246 1.475 0.279 ;
      RECT 1.426 0.175 1.437 0.304 ;
      RECT 0.993 0.246 1.126 0.279 ;
      RECT 2.547 0.17 3.022 0.26 ;
      RECT 1.437 0.17 2.044 0.26 ;
      RECT 0.635 0.17 1.031 0.26 ;
      RECT 1.38 0.204 2.044 0.26 ;
      RECT 1.464 1.14 2.119 1.23 ;
      RECT 2.029 0.85 2.119 1.23 ;
      RECT 2.549 1.092 2.779 1.182 ;
      RECT 2.54 1.049 2.549 1.178 ;
      RECT 2.54 1.092 2.825 1.159 ;
      RECT 2.502 1.092 2.825 1.154 ;
      RECT 1.464 0.525 1.554 1.23 ;
      RECT 2.029 1.045 2.54 1.135 ;
      RECT 0.148 1.045 1.554 1.135 ;
      RECT 2.741 1.073 2.871 1.113 ;
      RECT 2.029 1.073 2.587 1.135 ;
      RECT 2.779 1.031 2.871 1.113 ;
      RECT 0.148 0.943 0.238 1.135 ;
      RECT 0.045 0.943 0.238 1.033 ;
      RECT 2.825 0.985 2.918 1.044 ;
      RECT 2.871 0.939 2.917 1.067 ;
      RECT 2.825 0.985 2.956 1.024 ;
      RECT 3.252 0.702 3.342 1.005 ;
      RECT 2.917 0.915 3.342 1.005 ;
      RECT 0.045 0.335 0.135 1.033 ;
      RECT 1.979 0.85 2.119 0.94 ;
      RECT 1.464 0.525 1.654 0.665 ;
      RECT 0.455 0.476 0.545 0.66 ;
      RECT 0.428 0.394 0.455 0.523 ;
      RECT 0.382 0.358 0.428 0.486 ;
      RECT 0.382 0.431 0.501 0.486 ;
      RECT 0.344 0.335 0.382 0.444 ;
      RECT 0.045 0.335 0.382 0.425 ;
      RECT 1.669 0.96 1.834 1.05 ;
      RECT 1.744 0.35 1.834 1.05 ;
      RECT 2.444 0.67 2.534 0.821 ;
      RECT 1.744 0.67 2.534 0.76 ;
      RECT 1.694 0.35 1.834 0.44 ;
      RECT 0.884 0.865 1.364 0.955 ;
      RECT 1.274 0.621 1.364 0.955 ;
      RECT 1.188 0.621 1.364 0.711 ;
      RECT 1.144 0.561 1.188 0.689 ;
      RECT 1.098 0.516 1.144 0.644 ;
      RECT 1.098 0.602 1.226 0.644 ;
      RECT 1.052 0.47 1.098 0.598 ;
      RECT 1.006 0.424 1.052 0.552 ;
      RECT 0.96 0.378 1.006 0.506 ;
      RECT 0.922 0.424 1.052 0.464 ;
      RECT 0.82 0.355 0.96 0.445 ;
      RECT 3.541 0.17 4.667 0.26 ;
      RECT 4.037 0.9 4.457 0.99 ;
  END
END DFFRQX1H7R

MACRO DFFRQX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRQX2H7R 0 0 ;
  SIZE 5.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.6 1.48 ;
        RECT 5.415 1.225 5.555 1.48 ;
        RECT 4.527 1.225 4.667 1.48 ;
        RECT 2.864 1.225 3.004 1.48 ;
        RECT 2.324 1.225 2.464 1.48 ;
        RECT 1.164 1.225 1.304 1.48 ;
        RECT 0.31 1.225 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.6 0.08 ;
        RECT 5.072 -0.08 5.212 0.175 ;
        RECT 3.131 -0.08 3.271 0.175 ;
        RECT 2.299 -0.08 2.389 0.2 ;
        RECT 1.164 -0.08 1.304 0.175 ;
        RECT 0.31 -0.08 0.45 0.325 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.595 0.345 0.82 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.815 0.664 0.987 0.775 ;
        RECT 0.815 0.607 0.955 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.125 0.265 5.215 0.945 ;
        RECT 4.757 0.265 5.215 0.355 ;
        RECT 4.825 0.235 4.975 0.355 ;
      LAYER MET2 ;
        RECT 4.85 0.18 4.95 0.56 ;
      LAYER VIA1 ;
        RECT 4.855 0.255 4.945 0.345 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.995 0.625 3.145 0.805 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END RN
  OBS
    LAYER MET1 ;
      RECT 4.842 1.035 5.53 1.125 ;
      RECT 5.44 0.284 5.53 1.125 ;
      RECT 4.907 0.445 4.997 1.125 ;
      RECT 4.442 0.445 4.582 0.61 ;
      RECT 4.442 0.445 4.997 0.535 ;
      RECT 3.144 1.14 4.386 1.23 ;
      RECT 3.144 1.14 4.432 1.207 ;
      RECT 4.348 1.121 4.478 1.161 ;
      RECT 3.645 1.08 3.785 1.23 ;
      RECT 3.144 1.107 3.284 1.23 ;
      RECT 4.386 1.079 4.478 1.161 ;
      RECT 4.386 1.079 4.524 1.115 ;
      RECT 4.432 1.033 4.547 1.081 ;
      RECT 4.478 0.987 4.593 1.046 ;
      RECT 4.524 0.952 4.547 1.081 ;
      RECT 4.547 0.7 4.637 1.001 ;
      RECT 4.087 0.7 4.817 0.79 ;
      RECT 4.727 0.635 4.817 0.79 ;
      RECT 4.087 0.35 4.177 0.79 ;
      RECT 4.037 0.35 4.177 0.44 ;
      RECT 3.42 0.85 3.51 1.025 ;
      RECT 2.624 0.47 2.714 0.991 ;
      RECT 3.42 0.85 3.87 0.94 ;
      RECT 3.78 0.35 3.87 0.94 ;
      RECT 3.5 0.641 3.87 0.731 ;
      RECT 3.48 0.593 3.5 0.721 ;
      RECT 3.434 0.56 3.48 0.688 ;
      RECT 3.388 0.514 3.434 0.642 ;
      RECT 3.388 0.622 3.538 0.642 ;
      RECT 3.342 0.468 3.388 0.596 ;
      RECT 2.189 0.47 2.714 0.56 ;
      RECT 3.304 0.514 3.434 0.554 ;
      RECT 2.634 0.445 3.342 0.535 ;
      RECT 2.634 0.35 2.774 0.535 ;
      RECT 3.78 0.35 3.926 0.44 ;
      RECT 0.57 0.865 0.725 0.955 ;
      RECT 0.635 0.17 0.725 0.955 ;
      RECT 1.929 0.48 2.069 0.57 ;
      RECT 1.979 0.17 2.069 0.57 ;
      RECT 3.581 0.375 3.671 0.515 ;
      RECT 3.49 0.375 3.671 0.465 ;
      RECT 3.464 0.324 3.49 0.452 ;
      RECT 3.418 0.288 3.464 0.416 ;
      RECT 1.979 0.29 2.465 0.38 ;
      RECT 0.575 0.285 0.725 0.375 ;
      RECT 3.418 0.356 3.528 0.416 ;
      RECT 3.38 0.265 3.418 0.374 ;
      RECT 1.979 0.29 2.511 0.357 ;
      RECT 2.932 0.265 3.418 0.355 ;
      RECT 1.088 0.265 1.38 0.355 ;
      RECT 1.077 0.221 1.088 0.35 ;
      RECT 1.077 0.265 1.426 0.332 ;
      RECT 1.031 0.193 1.077 0.321 ;
      RECT 2.427 0.271 2.547 0.316 ;
      RECT 2.465 0.229 2.585 0.279 ;
      RECT 2.511 0.188 2.547 0.316 ;
      RECT 2.932 0.17 3.022 0.355 ;
      RECT 1.342 0.246 1.475 0.279 ;
      RECT 1.426 0.175 1.437 0.304 ;
      RECT 0.993 0.246 1.126 0.279 ;
      RECT 2.547 0.17 3.022 0.26 ;
      RECT 1.437 0.17 2.069 0.26 ;
      RECT 0.635 0.17 1.031 0.26 ;
      RECT 1.38 0.204 2.069 0.26 ;
      RECT 1.464 1.14 2.119 1.23 ;
      RECT 2.029 0.85 2.119 1.23 ;
      RECT 2.549 1.092 2.779 1.182 ;
      RECT 2.54 1.049 2.549 1.178 ;
      RECT 2.502 1.092 2.807 1.154 ;
      RECT 1.464 0.525 1.554 1.23 ;
      RECT 2.029 1.045 2.54 1.135 ;
      RECT 0.148 1.045 1.554 1.135 ;
      RECT 2.741 1.073 2.853 1.131 ;
      RECT 2.779 1.04 2.807 1.168 ;
      RECT 2.029 1.073 2.587 1.135 ;
      RECT 2.807 0.915 2.897 1.086 ;
      RECT 0.148 0.943 0.238 1.135 ;
      RECT 0.045 0.943 0.238 1.033 ;
      RECT 2.807 0.915 3.33 1.005 ;
      RECT 3.24 0.722 3.33 1.005 ;
      RECT 0.045 0.335 0.135 1.033 ;
      RECT 1.979 0.85 2.119 0.94 ;
      RECT 0.455 0.479 0.545 0.694 ;
      RECT 1.464 0.525 1.654 0.665 ;
      RECT 0.424 0.479 0.545 0.521 ;
      RECT 0.045 0.415 0.462 0.505 ;
      RECT 0.045 0.438 0.508 0.505 ;
      RECT 0.045 0.335 0.185 0.505 ;
      RECT 1.669 0.96 1.834 1.05 ;
      RECT 1.744 0.35 1.834 1.05 ;
      RECT 2.444 0.67 2.534 0.835 ;
      RECT 1.744 0.67 2.534 0.76 ;
      RECT 1.694 0.35 1.834 0.44 ;
      RECT 0.884 0.865 1.364 0.955 ;
      RECT 1.274 0.621 1.364 0.955 ;
      RECT 1.188 0.621 1.364 0.711 ;
      RECT 1.144 0.561 1.188 0.689 ;
      RECT 1.098 0.516 1.144 0.644 ;
      RECT 1.098 0.602 1.226 0.644 ;
      RECT 1.052 0.47 1.098 0.598 ;
      RECT 1.006 0.424 1.052 0.552 ;
      RECT 0.96 0.378 1.006 0.506 ;
      RECT 0.922 0.424 1.052 0.464 ;
      RECT 0.82 0.355 0.96 0.445 ;
      RECT 3.541 0.17 4.667 0.26 ;
      RECT 3.96 0.89 4.38 0.98 ;
  END
END DFFRQX2H7R

MACRO DFFRX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRX0P5H7R 0 0 ;
  SIZE 7 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7 1.48 ;
        RECT 6.495 1.195 6.635 1.48 ;
        RECT 5.71 1.225 5.85 1.48 ;
        RECT 4.452 1.225 4.592 1.48 ;
        RECT 2.225 0.89 2.315 1.48 ;
        RECT 0.805 1.225 0.945 1.48 ;
        RECT 0.335 1.165 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7 0.08 ;
        RECT 6.505 -0.08 6.595 0.385 ;
        RECT 6.015 -0.08 6.105 0.385 ;
        RECT 5.232 -0.08 5.375 0.175 ;
        RECT 4.462 -0.08 4.602 0.175 ;
        RECT 2.045 -0.08 2.135 0.385 ;
        RECT 0.845 -0.08 0.935 0.365 ;
        RECT 0.32 -0.08 0.41 0.335 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.35 0.695 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.73 1.175 0.945 ;
        RECT 0.92 0.685 1.115 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.792 0.425 6.945 0.575 ;
        RECT 6.792 0.31 6.882 0.925 ;
      LAYER MET2 ;
        RECT 6.85 0.23 6.95 0.76 ;
      LAYER VIA1 ;
        RECT 6.855 0.455 6.945 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.255 0.31 6.345 0.925 ;
      LAYER MET2 ;
        RECT 6.25 0.425 6.35 0.96 ;
      LAYER VIA1 ;
        RECT 6.255 0.655 6.345 0.745 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.705 0.455 3.795 0.865 ;
        RECT 3.625 0.455 3.795 0.545 ;
      LAYER MET2 ;
        RECT 3.65 0.23 3.75 0.76 ;
      LAYER VIA1 ;
        RECT 3.655 0.455 3.745 0.545 ;
    END
  END RN
  OBS
    LAYER MET1 ;
      RECT 6.015 1.015 6.68 1.105 ;
      RECT 6.59 0.575 6.68 1.105 ;
      RECT 6.015 0.626 6.105 1.105 ;
      RECT 5.993 0.547 6.015 0.675 ;
      RECT 5.947 0.513 5.993 0.641 ;
      RECT 5.947 0.581 6.061 0.641 ;
      RECT 5.901 0.467 5.947 0.595 ;
      RECT 5.855 0.421 5.901 0.549 ;
      RECT 5.811 0.17 5.855 0.504 ;
      RECT 5.765 0.17 5.855 0.459 ;
      RECT 5.555 0.17 5.855 0.26 ;
      RECT 5.082 1.045 5.172 1.23 ;
      RECT 5.082 1.045 5.855 1.135 ;
      RECT 5.765 0.655 5.855 1.135 ;
      RECT 3.445 0.78 3.59 0.87 ;
      RECT 3.445 0.17 3.535 0.87 ;
      RECT 5.376 0.655 5.855 0.745 ;
      RECT 5.376 0.305 5.466 0.745 ;
      RECT 4.423 0.305 5.466 0.395 ;
      RECT 4.418 0.264 4.423 0.393 ;
      RECT 4.372 0.239 4.418 0.367 ;
      RECT 4.326 0.193 4.372 0.321 ;
      RECT 4.326 0.286 4.461 0.321 ;
      RECT 4.288 0.17 4.326 0.279 ;
      RECT 3.445 0.17 4.326 0.26 ;
      RECT 2.855 0.96 4.236 1.05 ;
      RECT 2.855 0.96 4.282 1.027 ;
      RECT 4.198 0.941 4.331 0.974 ;
      RECT 4.282 0.87 4.293 0.999 ;
      RECT 2.855 0.93 2.995 1.05 ;
      RECT 5.532 0.835 5.672 0.955 ;
      RECT 4.236 0.899 5.672 0.955 ;
      RECT 4.293 0.865 5.672 0.955 ;
      RECT 4.262 0.665 5.282 0.755 ;
      RECT 4.255 0.623 4.262 0.752 ;
      RECT 4.217 0.665 5.282 0.729 ;
      RECT 4.107 0.62 4.255 0.71 ;
      RECT 4.107 0.646 4.3 0.71 ;
      RECT 2.44 1.14 4.316 1.23 ;
      RECT 2.44 1.14 4.362 1.207 ;
      RECT 4.882 1.045 4.972 1.195 ;
      RECT 4.278 1.121 4.411 1.154 ;
      RECT 4.362 1.05 4.373 1.179 ;
      RECT 4.373 1.045 4.972 1.135 ;
      RECT 4.316 1.079 4.972 1.135 ;
      RECT 3.91 0.78 4.05 0.87 ;
      RECT 3.91 0.476 4 0.87 ;
      RECT 4.347 0.485 4.691 0.575 ;
      RECT 4.306 0.426 4.347 0.555 ;
      RECT 3.91 0.476 4.046 0.514 ;
      RECT 4.26 0.383 4.306 0.511 ;
      RECT 4.26 0.466 4.385 0.511 ;
      RECT 3.956 0.431 4.049 0.49 ;
      RECT 4.222 0.36 4.26 0.469 ;
      RECT 3.956 0.431 4.087 0.469 ;
      RECT 4.049 0.36 4.26 0.45 ;
      RECT 4.046 0.361 4.049 0.49 ;
      RECT 4 0.386 4.306 0.45 ;
      RECT 3.14 0.78 3.285 0.87 ;
      RECT 3.195 0.255 3.285 0.87 ;
      RECT 2.42 0.495 3.285 0.585 ;
      RECT 2.42 0.32 2.51 0.585 ;
      RECT 2.27 0.32 2.51 0.41 ;
      RECT 1.035 1.14 2.135 1.23 ;
      RECT 2.045 0.7 2.135 1.23 ;
      RECT 1.035 1.045 1.125 1.23 ;
      RECT 0.956 1.045 1.125 1.135 ;
      RECT 0.938 0.998 0.956 1.126 ;
      RECT 0.892 0.966 0.938 1.094 ;
      RECT 0.846 0.92 0.892 1.048 ;
      RECT 0.846 1.026 0.994 1.048 ;
      RECT 0.8 0.874 0.846 1.002 ;
      RECT 0.754 0.828 0.8 0.956 ;
      RECT 0.716 0.874 0.846 0.914 ;
      RECT 0.5 0.805 0.754 0.895 ;
      RECT 2.96 0.675 3.05 0.815 ;
      RECT 0.5 0.285 0.59 0.895 ;
      RECT 2.045 0.7 3.05 0.79 ;
      RECT 0.5 0.285 0.715 0.375 ;
      RECT 2.63 0.88 2.72 1.05 ;
      RECT 2.405 0.88 2.72 0.97 ;
      RECT 1.435 0.935 1.955 1.025 ;
      RECT 1.865 0.52 1.955 1.025 ;
      RECT 1.435 0.35 1.525 1.025 ;
      RECT 1.865 0.52 2.27 0.61 ;
      RECT 1.385 0.35 1.525 0.44 ;
      RECT 1.685 0.17 1.775 0.83 ;
      RECT 1.205 0.17 1.295 0.64 ;
      RECT 0.69 0.505 1.295 0.595 ;
      RECT 1.205 0.17 1.775 0.26 ;
      RECT 0.515 1.12 0.655 1.21 ;
      RECT 0.515 0.985 0.605 1.21 ;
      RECT 0.07 0.985 0.605 1.075 ;
      RECT 0.07 0.26 0.16 1.075 ;
  END
END DFFRX0P5H7R

MACRO DFFRX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRX1H7R 0 0 ;
  SIZE 7 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7 1.48 ;
        RECT 6.5 1.195 6.64 1.48 ;
        RECT 5.71 1.225 5.85 1.48 ;
        RECT 4.452 1.225 4.592 1.48 ;
        RECT 2.225 0.89 2.315 1.48 ;
        RECT 0.805 1.225 0.945 1.48 ;
        RECT 0.335 1.165 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7 0.08 ;
        RECT 6.525 -0.08 6.615 0.345 ;
        RECT 6.015 -0.08 6.105 0.38 ;
        RECT 5.332 -0.08 5.422 0.345 ;
        RECT 4.462 -0.08 4.602 0.175 ;
        RECT 2.045 -0.08 2.135 0.38 ;
        RECT 0.845 -0.08 0.935 0.365 ;
        RECT 0.32 -0.08 0.41 0.335 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.35 0.695 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.73 1.175 0.945 ;
        RECT 0.92 0.685 1.115 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.792 0.425 6.945 0.575 ;
        RECT 6.792 0.31 6.882 0.925 ;
      LAYER MET2 ;
        RECT 6.85 0.23 6.95 0.76 ;
      LAYER VIA1 ;
        RECT 6.855 0.455 6.945 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.255 0.31 6.345 0.925 ;
      LAYER MET2 ;
        RECT 6.25 0.425 6.35 0.96 ;
      LAYER VIA1 ;
        RECT 6.255 0.655 6.345 0.745 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.705 0.455 3.795 0.865 ;
        RECT 3.625 0.455 3.795 0.545 ;
      LAYER MET2 ;
        RECT 3.65 0.23 3.75 0.76 ;
      LAYER VIA1 ;
        RECT 3.655 0.455 3.745 0.545 ;
    END
  END RN
  OBS
    LAYER MET1 ;
      RECT 6.015 1.015 6.68 1.105 ;
      RECT 6.59 0.575 6.68 1.105 ;
      RECT 6.015 0.576 6.105 1.105 ;
      RECT 5.972 0.486 6.015 0.615 ;
      RECT 5.972 0.531 6.061 0.615 ;
      RECT 5.926 0.442 5.972 0.57 ;
      RECT 5.88 0.396 5.926 0.524 ;
      RECT 5.866 0.305 5.88 0.494 ;
      RECT 5.82 0.305 5.88 0.464 ;
      RECT 5.774 0.305 5.88 0.418 ;
      RECT 5.54 0.305 5.88 0.395 ;
      RECT 5.057 1.045 5.91 1.135 ;
      RECT 5.82 0.639 5.91 1.135 ;
      RECT 3.445 0.78 3.59 0.87 ;
      RECT 3.445 0.17 3.535 0.87 ;
      RECT 5.78 0.551 5.82 0.679 ;
      RECT 5.78 0.594 5.866 0.679 ;
      RECT 5.734 0.508 5.78 0.636 ;
      RECT 5.696 0.485 5.734 0.594 ;
      RECT 5.101 0.485 5.734 0.575 ;
      RECT 5.101 0.265 5.191 0.575 ;
      RECT 4.383 0.265 5.191 0.355 ;
      RECT 4.372 0.221 4.383 0.35 ;
      RECT 4.326 0.193 4.372 0.321 ;
      RECT 4.777 0.24 4.917 0.355 ;
      RECT 4.288 0.246 4.421 0.279 ;
      RECT 3.445 0.17 4.326 0.26 ;
      RECT 2.855 0.96 4.141 1.05 ;
      RECT 2.855 0.96 4.187 1.027 ;
      RECT 4.103 0.941 4.236 0.974 ;
      RECT 4.187 0.87 4.198 0.999 ;
      RECT 2.855 0.93 2.995 1.05 ;
      RECT 5.532 0.835 5.672 0.955 ;
      RECT 4.141 0.899 5.672 0.955 ;
      RECT 4.198 0.865 5.672 0.955 ;
      RECT 4.262 0.665 5.282 0.755 ;
      RECT 4.255 0.623 4.262 0.752 ;
      RECT 4.217 0.665 5.282 0.729 ;
      RECT 4.107 0.62 4.255 0.71 ;
      RECT 4.107 0.646 4.3 0.71 ;
      RECT 2.44 1.14 4.236 1.23 ;
      RECT 2.44 1.14 4.282 1.207 ;
      RECT 4.872 1.045 4.962 1.195 ;
      RECT 4.198 1.121 4.331 1.154 ;
      RECT 4.282 1.05 4.293 1.179 ;
      RECT 4.293 1.045 4.962 1.135 ;
      RECT 4.236 1.079 4.962 1.135 ;
      RECT 3.91 0.78 4.05 0.87 ;
      RECT 3.91 0.476 4 0.87 ;
      RECT 4.345 0.485 4.741 0.575 ;
      RECT 4.304 0.426 4.345 0.555 ;
      RECT 3.91 0.476 4.046 0.514 ;
      RECT 4.258 0.383 4.304 0.511 ;
      RECT 4.258 0.466 4.383 0.511 ;
      RECT 3.956 0.431 4.049 0.49 ;
      RECT 4.22 0.36 4.258 0.469 ;
      RECT 3.956 0.431 4.087 0.469 ;
      RECT 4.049 0.36 4.258 0.45 ;
      RECT 4.046 0.361 4.049 0.49 ;
      RECT 4 0.386 4.304 0.45 ;
      RECT 3.14 0.78 3.285 0.87 ;
      RECT 3.195 0.275 3.285 0.87 ;
      RECT 2.415 0.495 3.285 0.585 ;
      RECT 2.415 0.32 2.505 0.585 ;
      RECT 2.27 0.32 2.505 0.41 ;
      RECT 1.035 1.14 2.135 1.23 ;
      RECT 2.045 0.7 2.135 1.23 ;
      RECT 1.035 1.045 1.125 1.23 ;
      RECT 0.921 1.045 1.125 1.135 ;
      RECT 0.903 0.998 0.921 1.126 ;
      RECT 0.857 0.966 0.903 1.094 ;
      RECT 0.811 0.92 0.857 1.048 ;
      RECT 0.811 1.026 0.959 1.048 ;
      RECT 0.765 0.874 0.811 1.002 ;
      RECT 0.719 0.828 0.765 0.956 ;
      RECT 0.681 0.874 0.811 0.914 ;
      RECT 0.5 0.805 0.719 0.895 ;
      RECT 2.96 0.675 3.05 0.815 ;
      RECT 0.5 0.285 0.59 0.895 ;
      RECT 2.045 0.7 3.05 0.79 ;
      RECT 0.5 0.285 0.715 0.375 ;
      RECT 2.63 0.88 2.72 1.045 ;
      RECT 2.405 0.88 2.72 0.97 ;
      RECT 1.435 0.935 1.955 1.025 ;
      RECT 1.865 0.52 1.955 1.025 ;
      RECT 1.435 0.35 1.525 1.025 ;
      RECT 1.865 0.52 2.27 0.61 ;
      RECT 1.385 0.35 1.525 0.44 ;
      RECT 1.685 0.17 1.775 0.83 ;
      RECT 1.205 0.17 1.295 0.64 ;
      RECT 0.69 0.5 1.295 0.59 ;
      RECT 1.205 0.17 1.775 0.26 ;
      RECT 0.515 1.12 0.655 1.21 ;
      RECT 0.515 0.985 0.605 1.21 ;
      RECT 0.07 0.985 0.605 1.075 ;
      RECT 0.07 0.26 0.16 1.075 ;
  END
END DFFRX1H7R

MACRO DFFRX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRX2H7R 0 0 ;
  SIZE 7.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7.4 1.48 ;
        RECT 7.22 1.035 7.31 1.48 ;
        RECT 6.68 1.225 6.82 1.48 ;
        RECT 5.82 1.225 5.96 1.48 ;
        RECT 4.597 1.225 4.737 1.48 ;
        RECT 2.37 0.89 2.46 1.48 ;
        RECT 0.975 1.2 1.065 1.48 ;
        RECT 0.335 1.175 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7.4 0.08 ;
        RECT 7.15 -0.08 7.24 0.33 ;
        RECT 6.64 -0.08 6.73 0.33 ;
        RECT 6.16 -0.08 6.25 0.36 ;
        RECT 5.407 -0.08 5.497 0.365 ;
        RECT 4.607 -0.08 4.752 0.175 ;
        RECT 2.12 -0.08 2.21 0.36 ;
        RECT 0.99 -0.08 1.08 0.345 ;
        RECT 0.32 -0.08 0.41 0.345 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.54 0.35 0.81 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.816 1.445 0.975 ;
        RECT 1.219 0.794 1.345 0.836 ;
        RECT 1.181 0.749 1.301 0.799 ;
        RECT 1.065 0.708 1.255 0.78 ;
        RECT 1.065 0.69 1.219 0.78 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.97 0.235 7.06 1.128 ;
        RECT 6.825 0.235 7.06 0.345 ;
      LAYER MET2 ;
        RECT 6.85 0.18 6.95 0.56 ;
      LAYER VIA1 ;
        RECT 6.855 0.255 6.945 0.345 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.365 0.855 6.575 0.95 ;
        RECT 6.39 0.335 6.48 0.95 ;
      LAYER MET2 ;
        RECT 6.45 0.625 6.55 1.16 ;
      LAYER VIA1 ;
        RECT 6.455 0.855 6.545 0.945 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.85 0.425 3.945 0.865 ;
      LAYER MET2 ;
        RECT 3.85 0.23 3.95 0.76 ;
      LAYER VIA1 ;
        RECT 3.855 0.455 3.945 0.545 ;
    END
  END RN
  OBS
    LAYER MET1 ;
      RECT 6.16 1.045 6.88 1.135 ;
      RECT 6.79 0.655 6.88 1.135 ;
      RECT 6.16 0.556 6.25 1.135 ;
      RECT 6.117 0.466 6.16 0.595 ;
      RECT 6.117 0.511 6.206 0.595 ;
      RECT 6.071 0.422 6.117 0.55 ;
      RECT 6.025 0.376 6.071 0.504 ;
      RECT 5.985 0.305 6.025 0.461 ;
      RECT 5.939 0.376 6.071 0.418 ;
      RECT 5.635 0.305 6.025 0.395 ;
      RECT 5.202 1.045 6.07 1.135 ;
      RECT 5.98 0.634 6.07 1.135 ;
      RECT 3.59 0.78 3.735 0.87 ;
      RECT 3.59 0.17 3.68 0.87 ;
      RECT 5.945 0.548 5.98 0.677 ;
      RECT 5.899 0.508 5.945 0.636 ;
      RECT 5.899 0.589 6.026 0.636 ;
      RECT 5.861 0.485 5.899 0.594 ;
      RECT 5.151 0.485 5.899 0.575 ;
      RECT 5.151 0.265 5.241 0.575 ;
      RECT 4.531 0.265 5.241 0.355 ;
      RECT 4.52 0.221 4.531 0.35 ;
      RECT 4.474 0.193 4.52 0.321 ;
      RECT 4.436 0.246 4.569 0.279 ;
      RECT 3.59 0.17 4.474 0.26 ;
      RECT 3 0.96 4.381 1.05 ;
      RECT 3 0.96 4.427 1.027 ;
      RECT 4.343 0.941 4.476 0.974 ;
      RECT 4.427 0.87 4.438 0.999 ;
      RECT 3 0.93 3.14 1.05 ;
      RECT 5.677 0.835 5.817 0.955 ;
      RECT 4.381 0.899 5.817 0.955 ;
      RECT 4.438 0.865 5.817 0.955 ;
      RECT 4.432 0.685 5.427 0.775 ;
      RECT 5.287 0.665 5.427 0.775 ;
      RECT 4.395 0.628 4.432 0.757 ;
      RECT 4.357 0.685 5.427 0.719 ;
      RECT 4.252 0.61 4.395 0.7 ;
      RECT 4.252 0.666 4.47 0.7 ;
      RECT 2.585 1.14 4.461 1.23 ;
      RECT 2.585 1.14 4.507 1.207 ;
      RECT 5.017 1.045 5.107 1.195 ;
      RECT 4.423 1.121 4.556 1.154 ;
      RECT 4.507 1.05 4.518 1.179 ;
      RECT 4.518 1.045 5.107 1.135 ;
      RECT 4.461 1.079 5.107 1.135 ;
      RECT 4.055 0.78 4.195 0.87 ;
      RECT 4.055 0.476 4.145 0.87 ;
      RECT 4.515 0.505 4.886 0.595 ;
      RECT 4.49 0.454 4.515 0.583 ;
      RECT 4.444 0.419 4.49 0.547 ;
      RECT 4.055 0.476 4.191 0.514 ;
      RECT 4.444 0.486 4.553 0.547 ;
      RECT 4.398 0.373 4.444 0.501 ;
      RECT 4.101 0.431 4.204 0.485 ;
      RECT 4.36 0.35 4.398 0.459 ;
      RECT 4.101 0.431 4.242 0.459 ;
      RECT 4.204 0.35 4.398 0.44 ;
      RECT 4.191 0.356 4.204 0.485 ;
      RECT 4.145 0.386 4.444 0.44 ;
      RECT 3.285 0.78 3.43 0.87 ;
      RECT 3.34 0.29 3.43 0.87 ;
      RECT 2.55 0.52 2.69 0.61 ;
      RECT 2.6 0.29 2.69 0.61 ;
      RECT 2.345 0.29 3.43 0.38 ;
      RECT 1.226 1.14 2.28 1.23 ;
      RECT 2.19 0.7 2.28 1.23 ;
      RECT 1.215 1.096 1.226 1.225 ;
      RECT 1.169 1.068 1.215 1.196 ;
      RECT 1.123 1.022 1.169 1.15 ;
      RECT 1.123 1.121 1.264 1.15 ;
      RECT 1.077 0.976 1.123 1.104 ;
      RECT 1.031 0.93 1.077 1.058 ;
      RECT 0.985 0.884 1.031 1.012 ;
      RECT 0.939 0.838 0.985 0.966 ;
      RECT 0.901 0.884 1.031 0.924 ;
      RECT 0.6 0.815 0.939 0.905 ;
      RECT 0.6 0.205 0.69 0.905 ;
      RECT 2.19 0.7 3.195 0.79 ;
      RECT 3.105 0.65 3.195 0.79 ;
      RECT 2.775 0.88 2.865 1.02 ;
      RECT 2.55 0.88 2.865 0.97 ;
      RECT 1.58 0.935 2.1 1.025 ;
      RECT 2.01 0.52 2.1 1.025 ;
      RECT 1.58 0.35 1.67 1.025 ;
      RECT 2.01 0.52 2.415 0.61 ;
      RECT 1.53 0.35 1.67 0.44 ;
      RECT 1.83 0.17 1.92 0.83 ;
      RECT 0.78 0.51 0.87 0.67 ;
      RECT 1.35 0.17 1.44 0.64 ;
      RECT 0.78 0.51 1.44 0.6 ;
      RECT 1.35 0.17 1.92 0.26 ;
      RECT 0.715 0.995 0.805 1.135 ;
      RECT 0.07 0.995 0.805 1.085 ;
      RECT 0.07 0.31 0.16 1.085 ;
  END
END DFFRX2H7R

MACRO DFFRX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRX3H7R 0 0 ;
  SIZE 7.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7.8 1.48 ;
        RECT 7.64 0.985 7.73 1.48 ;
        RECT 7.1 1.215 7.24 1.48 ;
        RECT 6.57 1.21 6.71 1.48 ;
        RECT 6.075 1.225 6.215 1.48 ;
        RECT 4.8 1.225 4.94 1.48 ;
        RECT 2.37 0.89 2.46 1.48 ;
        RECT 0.92 1.125 1.01 1.48 ;
        RECT 0.335 1.19 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7.8 0.08 ;
        RECT 7.64 -0.08 7.73 0.345 ;
        RECT 7.13 -0.08 7.22 0.33 ;
        RECT 6.63 -0.08 6.72 0.345 ;
        RECT 6.4 -0.08 6.49 0.345 ;
        RECT 5.725 -0.08 5.815 0.365 ;
        RECT 4.8 -0.08 4.94 0.175 ;
        RECT 2.12 -0.08 2.21 0.34 ;
        RECT 0.94 -0.08 1.03 0.345 ;
        RECT 0.32 -0.08 0.41 0.345 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.535 0.35 0.805 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.799 1.345 0.975 ;
        RECT 1.186 0.754 1.301 0.809 ;
        RECT 1.065 0.715 1.255 0.79 ;
        RECT 1.224 0.799 1.345 0.844 ;
        RECT 1.065 0.7 1.224 0.79 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.39 0.825 7.545 0.975 ;
        RECT 7.39 0.28 7.48 0.975 ;
      LAYER MET2 ;
        RECT 7.45 0.625 7.55 1.16 ;
      LAYER VIA1 ;
        RECT 7.455 0.855 7.545 0.945 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.825 0.855 6.975 0.945 ;
        RECT 6.88 0.28 6.975 0.945 ;
      LAYER MET2 ;
        RECT 6.85 0.63 6.95 1.16 ;
      LAYER VIA1 ;
        RECT 6.855 0.855 6.945 0.945 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.95 0.655 4.175 0.745 ;
        RECT 3.95 0.655 4.04 0.87 ;
      LAYER MET2 ;
        RECT 4.05 0.43 4.15 0.96 ;
      LAYER VIA1 ;
        RECT 4.055 0.655 4.145 0.745 ;
    END
  END RN
  OBS
    LAYER MET1 ;
      RECT 6.747 1.035 7.3 1.125 ;
      RECT 7.21 0.625 7.3 1.125 ;
      RECT 6.737 0.992 6.747 1.12 ;
      RECT 6.691 0.964 6.737 1.092 ;
      RECT 6.645 0.918 6.691 1.046 ;
      RECT 6.645 1.016 6.785 1.046 ;
      RECT 6.607 0.895 6.645 1.004 ;
      RECT 6.365 0.895 6.645 0.985 ;
      RECT 6.365 0.508 6.455 0.985 ;
      RECT 6.357 0.436 6.365 0.564 ;
      RECT 6.311 0.409 6.357 0.537 ;
      RECT 6.311 0.463 6.411 0.537 ;
      RECT 6.265 0.363 6.311 0.491 ;
      RECT 6.249 0.27 6.265 0.46 ;
      RECT 6.203 0.27 6.265 0.429 ;
      RECT 6.157 0.27 6.265 0.383 ;
      RECT 5.925 0.27 6.265 0.36 ;
      RECT 5.45 1.045 5.54 1.23 ;
      RECT 5.45 1.045 6.275 1.135 ;
      RECT 6.185 0.604 6.275 1.135 ;
      RECT 3.537 0.78 3.835 0.87 ;
      RECT 3.537 0.35 3.627 0.87 ;
      RECT 6.15 0.518 6.185 0.647 ;
      RECT 6.104 0.478 6.15 0.606 ;
      RECT 6.104 0.559 6.231 0.606 ;
      RECT 3.537 0.475 4.072 0.565 ;
      RECT 3.982 0.17 4.072 0.565 ;
      RECT 6.066 0.455 6.104 0.564 ;
      RECT 5.495 0.455 6.104 0.545 ;
      RECT 5.495 0.265 5.585 0.545 ;
      RECT 3.487 0.35 3.627 0.44 ;
      RECT 4.721 0.265 5.585 0.355 ;
      RECT 4.71 0.221 4.721 0.35 ;
      RECT 4.664 0.193 4.71 0.321 ;
      RECT 4.626 0.246 4.759 0.279 ;
      RECT 3.982 0.17 4.664 0.26 ;
      RECT 3 0.96 4.554 1.05 ;
      RECT 3 0.96 4.6 1.027 ;
      RECT 4.516 0.941 4.649 0.974 ;
      RECT 4.6 0.87 4.611 0.999 ;
      RECT 3 0.93 3.14 1.05 ;
      RECT 5.9 0.835 6.04 0.955 ;
      RECT 4.554 0.899 6.04 0.955 ;
      RECT 4.611 0.865 6.04 0.955 ;
      RECT 4.61 0.685 5.685 0.775 ;
      RECT 5.595 0.635 5.685 0.775 ;
      RECT 4.573 0.613 4.61 0.757 ;
      RECT 4.57 0.685 5.685 0.737 ;
      RECT 4.48 0.595 4.573 0.735 ;
      RECT 4.48 0.681 4.663 0.735 ;
      RECT 4.48 0.655 4.656 0.735 ;
      RECT 2.585 1.14 4.634 1.23 ;
      RECT 2.585 1.14 4.68 1.207 ;
      RECT 5.25 1.045 5.34 1.195 ;
      RECT 4.596 1.121 4.729 1.154 ;
      RECT 4.68 1.05 4.691 1.179 ;
      RECT 4.691 1.045 5.34 1.135 ;
      RECT 4.634 1.079 5.34 1.135 ;
      RECT 4.26 0.78 4.4 0.87 ;
      RECT 4.27 0.35 4.36 0.87 ;
      RECT 4.691 0.495 5.3 0.585 ;
      RECT 4.676 0.449 4.691 0.578 ;
      RECT 4.63 0.419 4.676 0.547 ;
      RECT 4.584 0.373 4.63 0.501 ;
      RECT 4.584 0.476 4.729 0.501 ;
      RECT 4.546 0.35 4.584 0.459 ;
      RECT 4.27 0.35 4.584 0.44 ;
      RECT 3.285 0.78 3.425 0.87 ;
      RECT 3.285 0.17 3.375 0.87 ;
      RECT 2.55 0.52 2.69 0.61 ;
      RECT 2.6 0.278 2.69 0.61 ;
      RECT 3.792 0.17 3.882 0.385 ;
      RECT 2.345 0.278 3.375 0.368 ;
      RECT 3.285 0.17 3.882 0.26 ;
      RECT 1.248 1.14 2.28 1.23 ;
      RECT 2.19 0.7 2.28 1.23 ;
      RECT 1.202 1.079 1.248 1.207 ;
      RECT 1.156 1.033 1.202 1.161 ;
      RECT 1.156 1.121 1.286 1.161 ;
      RECT 1.11 0.987 1.156 1.115 ;
      RECT 1.064 0.941 1.11 1.069 ;
      RECT 1.018 0.895 1.064 1.023 ;
      RECT 0.972 0.849 1.018 0.977 ;
      RECT 0.934 0.895 1.064 0.935 ;
      RECT 0.575 0.826 0.972 0.916 ;
      RECT 0.575 0.23 0.665 0.916 ;
      RECT 2.19 0.7 3.195 0.79 ;
      RECT 3.105 0.55 3.195 0.79 ;
      RECT 0.575 0.23 0.715 0.32 ;
      RECT 1.65 0.935 2.1 1.025 ;
      RECT 2.01 0.52 2.1 1.025 ;
      RECT 1.65 0.35 1.74 1.025 ;
      RECT 2.01 0.52 2.415 0.61 ;
      RECT 1.6 0.35 1.74 0.44 ;
      RECT 1.83 0.17 1.92 0.845 ;
      RECT 1.35 0.17 1.44 0.64 ;
      RECT 0.755 0.515 1.44 0.605 ;
      RECT 1.35 0.17 1.92 0.26 ;
      RECT 0.715 1.01 0.805 1.161 ;
      RECT 0.07 1.01 0.805 1.1 ;
      RECT 0.07 0.31 0.16 1.1 ;
      RECT 2.55 0.88 2.89 0.97 ;
  END
END DFFRX3H7R

MACRO DFFSQNX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSQNX1H7R 0 0 ;
  SIZE 5.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.8 1.48 ;
        RECT 5.315 1.225 5.455 1.48 ;
        RECT 4.785 1.225 4.925 1.48 ;
        RECT 4.164 1.225 4.304 1.48 ;
        RECT 1.953 1.225 2.093 1.48 ;
        RECT 0.815 1.225 0.955 1.48 ;
        RECT 0.31 1.225 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.8 0.08 ;
        RECT 5.246 -0.08 5.336 0.345 ;
        RECT 4.746 -0.08 4.836 0.33 ;
        RECT 3.916 -0.08 4.006 0.33 ;
        RECT 2.558 -0.08 2.698 0.175 ;
        RECT 1.95 -0.08 2.04 0.2 ;
        RECT 0.855 -0.08 0.945 0.345 ;
        RECT 0.352 -0.08 0.442 0.33 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.855 0.375 0.945 ;
        RECT 0.225 0.705 0.315 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.53 0.567 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.025 0.855 5.196 0.955 ;
        RECT 5.106 0.445 5.196 0.955 ;
        RECT 5.042 0.4 5.152 0.463 ;
        RECT 4.996 0.367 5.106 0.418 ;
        RECT 5.086 0.445 5.196 0.495 ;
        RECT 4.996 0.205 5.086 0.418 ;
      LAYER MET2 ;
        RECT 5.05 0.63 5.15 1.16 ;
      LAYER VIA1 ;
        RECT 5.055 0.855 5.145 0.945 ;
    END
  END QN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.445 0.425 5.545 0.695 ;
      LAYER MET2 ;
        RECT 5.45 0.225 5.55 0.76 ;
      LAYER VIA1 ;
        RECT 5.455 0.455 5.545 0.545 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 4.334 1.045 5.385 1.135 ;
      RECT 5.295 0.88 5.385 1.135 ;
      RECT 5.295 0.88 5.725 0.97 ;
      RECT 5.635 0.23 5.725 0.97 ;
      RECT 5.519 0.23 5.725 0.32 ;
      RECT 3.791 1.14 4.03 1.23 ;
      RECT 3.791 1.14 4.076 1.207 ;
      RECT 3.992 1.121 4.122 1.161 ;
      RECT 4.03 1.079 4.141 1.129 ;
      RECT 4.076 1.033 4.187 1.096 ;
      RECT 4.122 1 4.141 1.129 ;
      RECT 4.141 0.865 4.231 1.051 ;
      RECT 4.141 0.865 4.656 0.955 ;
      RECT 4.566 0.23 4.656 0.955 ;
      RECT 4.566 0.655 4.986 0.745 ;
      RECT 4.896 0.605 4.986 0.745 ;
      RECT 4.471 0.23 4.656 0.32 ;
      RECT 3.431 0.805 3.521 1.012 ;
      RECT 3.477 0.76 3.567 0.843 ;
      RECT 3.521 0.715 3.613 0.797 ;
      RECT 3.521 0.715 3.659 0.751 ;
      RECT 3.567 0.669 3.676 0.72 ;
      RECT 3.613 0.623 3.722 0.688 ;
      RECT 3.659 0.591 3.676 0.72 ;
      RECT 3.613 0.623 3.748 0.652 ;
      RECT 3.676 0.549 4.476 0.639 ;
      RECT 4.174 0.205 4.264 0.639 ;
      RECT 3.676 0.219 3.766 0.639 ;
      RECT 3.319 0.219 3.766 0.309 ;
      RECT 2.765 1.14 3.701 1.23 ;
      RECT 2.758 1.098 2.765 1.227 ;
      RECT 2.72 1.14 3.701 1.204 ;
      RECT 2.618 1.095 2.758 1.185 ;
      RECT 3.611 0.975 3.701 1.23 ;
      RECT 2.618 1.121 2.803 1.185 ;
      RECT 3.611 0.975 3.753 1.003 ;
      RECT 3.715 0.894 4.006 0.984 ;
      RECT 3.657 0.93 4.006 0.984 ;
      RECT 3.701 0.901 3.715 1.029 ;
      RECT 2.183 1.045 2.323 1.23 ;
      RECT 1.195 1.14 1.755 1.23 ;
      RECT 1.665 1.045 1.755 1.23 ;
      RECT 1.195 0.475 1.285 1.23 ;
      RECT 1.665 1.045 2.44 1.135 ;
      RECT 0.045 1.045 1.285 1.135 ;
      RECT 1.665 1.045 2.496 1.102 ;
      RECT 2.45 0.83 2.54 1.057 ;
      RECT 2.841 0.96 3.311 1.05 ;
      RECT 2.402 1.026 2.54 1.057 ;
      RECT 2.44 1.002 2.45 1.13 ;
      RECT 0.045 0.246 0.135 1.135 ;
      RECT 2.795 0.899 2.841 1.027 ;
      RECT 2.749 0.853 2.795 0.981 ;
      RECT 3.221 0.759 3.311 1.05 ;
      RECT 2.749 0.941 2.879 0.981 ;
      RECT 2.711 0.899 2.841 0.939 ;
      RECT 2.45 0.83 2.749 0.92 ;
      RECT 3.221 0.759 3.357 0.797 ;
      RECT 3.267 0.714 3.374 0.766 ;
      RECT 3.311 0.669 3.42 0.734 ;
      RECT 3.357 0.637 3.374 0.766 ;
      RECT 3.374 0.419 3.464 0.689 ;
      RECT 3.374 0.419 3.529 0.509 ;
      RECT 0.045 0.246 0.217 0.336 ;
      RECT 1.555 0.865 2.358 0.955 ;
      RECT 1.555 0.47 1.645 0.955 ;
      RECT 1.555 0.47 2.34 0.56 ;
      RECT 2.249 0.375 2.34 0.56 ;
      RECT 3.139 0.17 3.229 0.555 ;
      RECT 2.249 0.375 2.664 0.465 ;
      RECT 2.249 0.375 2.71 0.442 ;
      RECT 2.626 0.356 2.756 0.396 ;
      RECT 2.664 0.314 2.756 0.396 ;
      RECT 2.71 0.268 2.802 0.35 ;
      RECT 2.756 0.222 2.869 0.279 ;
      RECT 2.802 0.184 2.831 0.313 ;
      RECT 2.831 0.17 3.229 0.26 ;
      RECT 2.937 0.78 3.077 0.87 ;
      RECT 2.937 0.35 3.027 0.87 ;
      RECT 1.819 0.65 3.027 0.74 ;
      RECT 2.909 0.35 3.049 0.44 ;
      RECT 1.375 0.22 1.465 1.02 ;
      RECT 1.375 0.29 2.116 0.38 ;
      RECT 1.375 0.29 2.162 0.357 ;
      RECT 2.078 0.271 2.198 0.316 ;
      RECT 2.116 0.229 2.236 0.279 ;
      RECT 2.162 0.188 2.198 0.316 ;
      RECT 2.198 0.17 2.468 0.26 ;
      RECT 0.625 0.865 0.765 0.955 ;
      RECT 0.657 0.651 0.765 0.955 ;
      RECT 0.657 0.651 1.05 0.741 ;
      RECT 0.657 0.29 0.747 0.955 ;
      RECT 0.599 0.29 0.747 0.38 ;
  END
END DFFSQNX1H7R

MACRO DFFSQNX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSQNX2H7R 0 0 ;
  SIZE 5.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.8 1.48 ;
        RECT 5.315 1.225 5.455 1.48 ;
        RECT 4.785 1.225 4.925 1.48 ;
        RECT 4.164 1.225 4.304 1.48 ;
        RECT 1.953 1.225 2.093 1.48 ;
        RECT 0.815 1.225 0.955 1.48 ;
        RECT 0.31 1.225 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.8 0.08 ;
        RECT 5.246 -0.08 5.336 0.33 ;
        RECT 4.746 -0.08 4.836 0.33 ;
        RECT 3.916 -0.08 4.006 0.33 ;
        RECT 2.558 -0.08 2.698 0.175 ;
        RECT 1.95 -0.08 2.04 0.2 ;
        RECT 0.855 -0.08 0.945 0.345 ;
        RECT 0.352 -0.08 0.442 0.33 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.855 0.375 0.945 ;
        RECT 0.225 0.705 0.315 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.53 0.567 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.025 0.855 5.196 0.955 ;
        RECT 5.106 0.445 5.196 0.955 ;
        RECT 5.042 0.4 5.152 0.463 ;
        RECT 4.996 0.367 5.106 0.418 ;
        RECT 5.086 0.445 5.196 0.495 ;
        RECT 4.996 0.22 5.086 0.418 ;
      LAYER MET2 ;
        RECT 5.05 0.63 5.15 1.16 ;
      LAYER VIA1 ;
        RECT 5.055 0.855 5.145 0.945 ;
    END
  END QN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.445 0.425 5.545 0.695 ;
      LAYER MET2 ;
        RECT 5.45 0.225 5.55 0.76 ;
      LAYER VIA1 ;
        RECT 5.455 0.455 5.545 0.545 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 4.334 1.045 5.385 1.135 ;
      RECT 5.295 0.88 5.385 1.135 ;
      RECT 5.295 0.88 5.725 0.97 ;
      RECT 5.635 0.23 5.725 0.97 ;
      RECT 5.519 0.23 5.725 0.32 ;
      RECT 3.791 1.14 4.03 1.23 ;
      RECT 3.791 1.14 4.076 1.207 ;
      RECT 3.992 1.121 4.122 1.161 ;
      RECT 4.03 1.079 4.141 1.129 ;
      RECT 4.076 1.033 4.187 1.096 ;
      RECT 4.122 1 4.141 1.129 ;
      RECT 4.141 0.865 4.231 1.051 ;
      RECT 4.141 0.865 4.656 0.955 ;
      RECT 4.566 0.25 4.656 0.955 ;
      RECT 4.566 0.655 5.016 0.745 ;
      RECT 4.926 0.605 5.016 0.745 ;
      RECT 4.471 0.25 4.656 0.34 ;
      RECT 3.431 0.805 3.521 1.012 ;
      RECT 3.477 0.76 3.567 0.843 ;
      RECT 3.521 0.715 3.613 0.797 ;
      RECT 3.521 0.715 3.659 0.751 ;
      RECT 3.567 0.669 3.676 0.72 ;
      RECT 3.613 0.623 3.722 0.688 ;
      RECT 3.659 0.591 3.676 0.72 ;
      RECT 3.613 0.623 3.748 0.652 ;
      RECT 3.676 0.549 4.476 0.639 ;
      RECT 4.174 0.245 4.264 0.639 ;
      RECT 3.676 0.219 3.766 0.639 ;
      RECT 3.319 0.219 3.766 0.309 ;
      RECT 2.765 1.14 3.701 1.23 ;
      RECT 2.758 1.098 2.765 1.227 ;
      RECT 2.72 1.14 3.701 1.204 ;
      RECT 2.618 1.095 2.758 1.185 ;
      RECT 3.611 0.975 3.701 1.23 ;
      RECT 2.618 1.121 2.803 1.185 ;
      RECT 3.611 0.975 3.753 1.003 ;
      RECT 3.715 0.894 4.006 0.984 ;
      RECT 3.657 0.93 4.006 0.984 ;
      RECT 3.701 0.901 3.715 1.029 ;
      RECT 2.183 1.045 2.323 1.23 ;
      RECT 1.195 1.14 1.755 1.23 ;
      RECT 1.665 1.045 1.755 1.23 ;
      RECT 1.195 0.475 1.285 1.23 ;
      RECT 1.665 1.045 2.44 1.135 ;
      RECT 0.045 1.045 1.285 1.135 ;
      RECT 1.665 1.045 2.496 1.102 ;
      RECT 2.45 0.83 2.54 1.057 ;
      RECT 2.841 0.96 3.311 1.05 ;
      RECT 2.402 1.026 2.54 1.057 ;
      RECT 2.44 1.002 2.45 1.13 ;
      RECT 0.045 0.246 0.135 1.135 ;
      RECT 2.795 0.899 2.841 1.027 ;
      RECT 2.749 0.853 2.795 0.981 ;
      RECT 3.221 0.759 3.311 1.05 ;
      RECT 2.749 0.941 2.879 0.981 ;
      RECT 2.711 0.899 2.841 0.939 ;
      RECT 2.45 0.83 2.749 0.92 ;
      RECT 3.221 0.759 3.357 0.797 ;
      RECT 3.267 0.714 3.374 0.766 ;
      RECT 3.311 0.669 3.42 0.734 ;
      RECT 3.357 0.637 3.374 0.766 ;
      RECT 3.374 0.419 3.464 0.689 ;
      RECT 3.374 0.419 3.529 0.509 ;
      RECT 0.045 0.246 0.217 0.336 ;
      RECT 1.555 0.865 2.358 0.955 ;
      RECT 1.555 0.47 1.645 0.955 ;
      RECT 1.555 0.47 2.34 0.56 ;
      RECT 2.249 0.375 2.34 0.56 ;
      RECT 3.139 0.17 3.229 0.555 ;
      RECT 2.249 0.375 2.664 0.465 ;
      RECT 2.249 0.375 2.71 0.442 ;
      RECT 2.626 0.356 2.756 0.396 ;
      RECT 2.664 0.314 2.756 0.396 ;
      RECT 2.71 0.268 2.802 0.35 ;
      RECT 2.756 0.222 2.869 0.279 ;
      RECT 2.802 0.184 2.831 0.313 ;
      RECT 2.831 0.17 3.229 0.26 ;
      RECT 2.937 0.78 3.077 0.87 ;
      RECT 2.937 0.35 3.027 0.87 ;
      RECT 1.819 0.65 3.027 0.74 ;
      RECT 2.909 0.35 3.049 0.44 ;
      RECT 1.375 0.22 1.465 1.01 ;
      RECT 1.375 0.29 2.116 0.38 ;
      RECT 1.375 0.29 2.162 0.357 ;
      RECT 2.078 0.271 2.198 0.316 ;
      RECT 2.116 0.229 2.236 0.279 ;
      RECT 2.162 0.188 2.198 0.316 ;
      RECT 2.198 0.17 2.468 0.26 ;
      RECT 0.625 0.85 0.765 0.94 ;
      RECT 0.657 0.651 0.765 0.94 ;
      RECT 0.657 0.651 1.05 0.741 ;
      RECT 0.657 0.354 0.747 0.94 ;
      RECT 0.599 0.354 0.747 0.444 ;
  END
END DFFSQNX2H7R

MACRO DFFSQX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSQX1H7R 0 0 ;
  SIZE 5.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.8 1.48 ;
        RECT 5.315 1.225 5.455 1.48 ;
        RECT 4.785 1.225 4.925 1.48 ;
        RECT 4.164 1.225 4.304 1.48 ;
        RECT 1.953 1.225 2.093 1.48 ;
        RECT 0.815 1.225 0.955 1.48 ;
        RECT 0.31 1.225 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.8 0.08 ;
        RECT 5.246 -0.08 5.336 0.345 ;
        RECT 4.746 -0.08 4.836 0.33 ;
        RECT 3.916 -0.08 4.006 0.33 ;
        RECT 2.558 -0.08 2.698 0.175 ;
        RECT 1.95 -0.08 2.04 0.2 ;
        RECT 0.855 -0.08 0.945 0.345 ;
        RECT 0.352 -0.08 0.442 0.33 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.855 0.41 0.945 ;
        RECT 0.225 0.74 0.315 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.53 0.567 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.996 0.855 5.19 0.955 ;
        RECT 4.996 0.265 5.086 0.955 ;
      LAYER MET2 ;
        RECT 5.05 0.63 5.15 1.16 ;
      LAYER VIA1 ;
        RECT 5.055 0.855 5.145 0.945 ;
    END
  END Q
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.365 0.625 5.545 0.775 ;
      LAYER MET2 ;
        RECT 5.45 0.425 5.55 0.96 ;
      LAYER VIA1 ;
        RECT 5.455 0.655 5.545 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 4.334 1.045 5.37 1.135 ;
      RECT 5.28 0.88 5.37 1.135 ;
      RECT 5.28 0.88 5.725 0.97 ;
      RECT 5.635 0.23 5.725 0.97 ;
      RECT 5.519 0.23 5.725 0.32 ;
      RECT 3.791 1.14 4.03 1.23 ;
      RECT 3.791 1.14 4.076 1.207 ;
      RECT 3.992 1.121 4.122 1.161 ;
      RECT 4.03 1.079 4.141 1.129 ;
      RECT 4.076 1.033 4.187 1.096 ;
      RECT 4.122 1 4.141 1.129 ;
      RECT 4.141 0.865 4.231 1.051 ;
      RECT 4.141 0.865 4.656 0.955 ;
      RECT 4.566 0.23 4.656 0.955 ;
      RECT 4.471 0.23 4.656 0.32 ;
      RECT 3.431 0.805 3.521 1.012 ;
      RECT 3.477 0.76 3.567 0.843 ;
      RECT 3.521 0.715 3.613 0.797 ;
      RECT 3.521 0.715 3.659 0.751 ;
      RECT 3.567 0.669 3.676 0.72 ;
      RECT 3.613 0.623 3.722 0.688 ;
      RECT 3.659 0.591 3.676 0.72 ;
      RECT 3.613 0.623 3.748 0.652 ;
      RECT 3.676 0.549 4.476 0.639 ;
      RECT 4.174 0.205 4.264 0.639 ;
      RECT 3.676 0.219 3.766 0.639 ;
      RECT 3.319 0.219 3.766 0.309 ;
      RECT 2.765 1.14 3.701 1.23 ;
      RECT 2.758 1.098 2.765 1.227 ;
      RECT 2.72 1.14 3.701 1.204 ;
      RECT 2.618 1.095 2.758 1.185 ;
      RECT 3.611 0.975 3.701 1.23 ;
      RECT 2.618 1.121 2.803 1.185 ;
      RECT 3.611 0.975 3.753 1.003 ;
      RECT 3.715 0.894 4.006 0.984 ;
      RECT 3.657 0.93 4.006 0.984 ;
      RECT 3.701 0.901 3.715 1.029 ;
      RECT 2.183 1.045 2.323 1.23 ;
      RECT 1.12 1.14 1.755 1.23 ;
      RECT 1.665 1.045 1.755 1.23 ;
      RECT 1.12 0.658 1.21 1.23 ;
      RECT 1.665 1.045 2.44 1.135 ;
      RECT 0.045 1.045 1.21 1.135 ;
      RECT 1.665 1.045 2.496 1.102 ;
      RECT 2.45 0.83 2.54 1.057 ;
      RECT 2.841 0.96 3.311 1.05 ;
      RECT 2.402 1.026 2.54 1.057 ;
      RECT 2.44 1.002 2.45 1.13 ;
      RECT 0.045 0.246 0.135 1.135 ;
      RECT 2.795 0.899 2.841 1.027 ;
      RECT 2.749 0.853 2.795 0.981 ;
      RECT 3.221 0.759 3.311 1.05 ;
      RECT 2.749 0.941 2.879 0.981 ;
      RECT 2.711 0.899 2.841 0.939 ;
      RECT 2.45 0.83 2.749 0.92 ;
      RECT 3.221 0.759 3.357 0.797 ;
      RECT 3.267 0.714 3.374 0.766 ;
      RECT 1.195 0.475 1.285 0.748 ;
      RECT 3.311 0.669 3.42 0.734 ;
      RECT 3.357 0.637 3.374 0.766 ;
      RECT 3.374 0.419 3.464 0.689 ;
      RECT 3.374 0.419 3.529 0.509 ;
      RECT 0.045 0.246 0.217 0.336 ;
      RECT 1.555 0.865 2.358 0.955 ;
      RECT 1.555 0.47 1.645 0.955 ;
      RECT 1.555 0.47 2.339 0.56 ;
      RECT 2.249 0.375 2.339 0.56 ;
      RECT 3.139 0.17 3.229 0.555 ;
      RECT 2.249 0.375 2.664 0.465 ;
      RECT 2.249 0.375 2.71 0.442 ;
      RECT 2.626 0.356 2.756 0.396 ;
      RECT 2.664 0.314 2.756 0.396 ;
      RECT 2.71 0.268 2.802 0.35 ;
      RECT 2.756 0.222 2.869 0.279 ;
      RECT 2.802 0.184 2.831 0.313 ;
      RECT 2.831 0.17 3.229 0.26 ;
      RECT 2.937 0.78 3.077 0.87 ;
      RECT 2.937 0.35 3.027 0.87 ;
      RECT 1.819 0.65 3.027 0.74 ;
      RECT 2.909 0.35 3.049 0.44 ;
      RECT 1.3 0.89 1.465 0.98 ;
      RECT 1.375 0.22 1.465 0.98 ;
      RECT 1.375 0.29 2.116 0.38 ;
      RECT 1.375 0.29 2.162 0.357 ;
      RECT 2.078 0.271 2.198 0.316 ;
      RECT 2.116 0.229 2.236 0.279 ;
      RECT 2.162 0.188 2.198 0.316 ;
      RECT 2.198 0.17 2.468 0.26 ;
      RECT 0.625 0.865 0.765 0.955 ;
      RECT 0.657 0.651 0.765 0.955 ;
      RECT 0.657 0.651 1.01 0.741 ;
      RECT 0.657 0.29 0.747 0.955 ;
      RECT 0.599 0.29 0.747 0.38 ;
  END
END DFFSQX1H7R

MACRO DFFSQX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSQX2H7R 0 0 ;
  SIZE 5.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.8 1.48 ;
        RECT 5.315 1.225 5.455 1.48 ;
        RECT 4.785 1.225 4.925 1.48 ;
        RECT 4.164 1.225 4.304 1.48 ;
        RECT 1.934 1.225 2.093 1.48 ;
        RECT 0.815 1.225 0.955 1.48 ;
        RECT 0.31 1.225 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.8 0.08 ;
        RECT 5.246 -0.08 5.336 0.33 ;
        RECT 4.746 -0.08 4.836 0.33 ;
        RECT 3.916 -0.08 4.006 0.33 ;
        RECT 2.558 -0.08 2.698 0.175 ;
        RECT 1.95 -0.08 2.04 0.2 ;
        RECT 0.855 -0.08 0.945 0.345 ;
        RECT 0.352 -0.08 0.442 0.33 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.855 0.41 0.945 ;
        RECT 0.225 0.74 0.315 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.53 0.567 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.996 0.855 5.19 0.955 ;
        RECT 4.996 0.22 5.086 0.955 ;
      LAYER MET2 ;
        RECT 5.05 0.63 5.15 1.16 ;
      LAYER VIA1 ;
        RECT 5.055 0.855 5.145 0.945 ;
    END
  END Q
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.365 0.625 5.545 0.775 ;
      LAYER MET2 ;
        RECT 5.45 0.425 5.55 0.96 ;
      LAYER VIA1 ;
        RECT 5.455 0.655 5.545 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 4.334 1.045 5.37 1.135 ;
      RECT 5.28 0.88 5.37 1.135 ;
      RECT 5.28 0.88 5.725 0.97 ;
      RECT 5.635 0.23 5.725 0.97 ;
      RECT 5.519 0.23 5.725 0.32 ;
      RECT 3.791 1.14 4.03 1.23 ;
      RECT 3.791 1.14 4.076 1.207 ;
      RECT 3.992 1.121 4.122 1.161 ;
      RECT 4.03 1.079 4.141 1.129 ;
      RECT 4.076 1.033 4.187 1.096 ;
      RECT 4.122 1 4.141 1.129 ;
      RECT 4.141 0.865 4.231 1.051 ;
      RECT 4.141 0.865 4.656 0.955 ;
      RECT 4.566 0.25 4.656 0.955 ;
      RECT 4.471 0.25 4.656 0.34 ;
      RECT 3.431 0.805 3.521 1.012 ;
      RECT 3.477 0.76 3.567 0.843 ;
      RECT 3.521 0.715 3.613 0.797 ;
      RECT 3.521 0.715 3.659 0.751 ;
      RECT 3.567 0.669 3.676 0.72 ;
      RECT 3.613 0.623 3.722 0.688 ;
      RECT 3.659 0.591 3.676 0.72 ;
      RECT 3.613 0.623 3.748 0.652 ;
      RECT 3.676 0.549 4.476 0.639 ;
      RECT 4.174 0.245 4.264 0.639 ;
      RECT 3.676 0.219 3.766 0.639 ;
      RECT 3.319 0.219 3.766 0.309 ;
      RECT 2.765 1.14 3.701 1.23 ;
      RECT 2.758 1.098 2.765 1.227 ;
      RECT 2.72 1.14 3.701 1.204 ;
      RECT 2.618 1.095 2.758 1.185 ;
      RECT 3.611 0.975 3.701 1.23 ;
      RECT 2.618 1.121 2.803 1.185 ;
      RECT 3.611 0.975 3.753 1.003 ;
      RECT 3.715 0.894 4.006 0.984 ;
      RECT 3.657 0.93 4.006 0.984 ;
      RECT 3.701 0.901 3.715 1.029 ;
      RECT 2.183 1.045 2.323 1.23 ;
      RECT 1.1 1.14 1.755 1.23 ;
      RECT 1.665 1.045 1.755 1.23 ;
      RECT 1.1 0.658 1.19 1.23 ;
      RECT 1.665 1.045 2.44 1.135 ;
      RECT 0.045 1.045 1.19 1.135 ;
      RECT 1.665 1.045 2.496 1.102 ;
      RECT 2.45 0.83 2.54 1.057 ;
      RECT 2.841 0.96 3.311 1.05 ;
      RECT 2.402 1.026 2.54 1.057 ;
      RECT 2.44 1.002 2.45 1.13 ;
      RECT 0.045 0.246 0.135 1.135 ;
      RECT 2.795 0.899 2.841 1.027 ;
      RECT 2.749 0.853 2.795 0.981 ;
      RECT 3.221 0.759 3.311 1.05 ;
      RECT 2.749 0.941 2.879 0.981 ;
      RECT 2.711 0.899 2.841 0.939 ;
      RECT 2.45 0.83 2.749 0.92 ;
      RECT 3.221 0.759 3.357 0.797 ;
      RECT 3.267 0.714 3.374 0.766 ;
      RECT 1.1 0.658 1.285 0.748 ;
      RECT 1.195 0.475 1.285 0.748 ;
      RECT 3.311 0.669 3.42 0.734 ;
      RECT 3.357 0.637 3.374 0.766 ;
      RECT 3.374 0.419 3.464 0.689 ;
      RECT 3.374 0.419 3.529 0.509 ;
      RECT 0.045 0.246 0.217 0.336 ;
      RECT 1.555 0.865 2.358 0.955 ;
      RECT 1.555 0.47 1.645 0.955 ;
      RECT 1.555 0.47 2.339 0.56 ;
      RECT 2.249 0.375 2.339 0.56 ;
      RECT 3.139 0.17 3.229 0.555 ;
      RECT 2.249 0.375 2.664 0.465 ;
      RECT 2.249 0.375 2.71 0.442 ;
      RECT 2.626 0.356 2.756 0.396 ;
      RECT 2.664 0.314 2.756 0.396 ;
      RECT 2.71 0.268 2.802 0.35 ;
      RECT 2.756 0.222 2.869 0.279 ;
      RECT 2.802 0.184 2.831 0.313 ;
      RECT 2.831 0.17 3.229 0.26 ;
      RECT 2.937 0.78 3.077 0.87 ;
      RECT 2.937 0.35 3.027 0.87 ;
      RECT 1.819 0.65 3.027 0.74 ;
      RECT 2.909 0.35 3.049 0.44 ;
      RECT 1.3 0.946 1.465 1.036 ;
      RECT 1.375 0.22 1.465 1.036 ;
      RECT 1.375 0.29 2.116 0.38 ;
      RECT 1.375 0.29 2.162 0.357 ;
      RECT 2.078 0.271 2.198 0.316 ;
      RECT 2.116 0.229 2.236 0.279 ;
      RECT 2.162 0.188 2.198 0.316 ;
      RECT 2.198 0.17 2.468 0.26 ;
      RECT 0.625 0.85 0.765 0.94 ;
      RECT 0.675 0.344 0.765 0.94 ;
      RECT 0.675 0.651 1.01 0.741 ;
      RECT 0.599 0.344 0.765 0.434 ;
  END
END DFFSQX2H7R

MACRO DFFSRQX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRQX1H7R 0 0 ;
  SIZE 6.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.6 1.48 ;
        RECT 6.148 1.095 6.288 1.48 ;
        RECT 5.344 1.24 5.484 1.48 ;
        RECT 4.354 1.24 4.494 1.48 ;
        RECT 1.465 1.24 1.605 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.6 0.08 ;
        RECT 6.148 -0.08 6.288 0.305 ;
        RECT 4.895 -0.08 5.035 0.175 ;
        RECT 1.455 -0.08 1.545 0.315 ;
        RECT 0.31 -0.08 0.45 0.193 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.66 0.25 1.975 0.345 ;
      LAYER MET2 ;
        RECT 1.85 0.18 1.95 0.56 ;
      LAYER VIA1 ;
        RECT 1.855 0.255 1.945 0.345 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.655 0.585 0.825 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.434 0.225 6.545 1.077 ;
      LAYER MET2 ;
        RECT 6.45 0.18 6.55 0.56 ;
      LAYER VIA1 ;
        RECT 6.455 0.255 6.545 0.345 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.15 0.625 5.375 0.766 ;
      LAYER MET2 ;
        RECT 5.25 0.425 5.35 0.96 ;
      LAYER VIA1 ;
        RECT 5.255 0.655 5.345 0.745 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.561 0.455 5.775 0.627 ;
      LAYER MET2 ;
        RECT 5.65 0.225 5.75 0.76 ;
      LAYER VIA1 ;
        RECT 5.655 0.455 5.745 0.545 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 4.614 1.14 5.226 1.23 ;
      RECT 3.887 1.14 4.235 1.23 ;
      RECT 4.572 1.14 5.268 1.209 ;
      RECT 3.887 1.14 4.277 1.209 ;
      RECT 4.534 1.14 5.306 1.169 ;
      RECT 3.887 1.14 4.315 1.169 ;
      RECT 5.188 1.121 6.038 1.15 ;
      RECT 4.197 1.121 4.652 1.15 ;
      RECT 5.226 1.081 6.038 1.15 ;
      RECT 4.235 1.081 4.614 1.15 ;
      RECT 5.268 1.06 6.038 1.15 ;
      RECT 4.277 1.06 4.572 1.15 ;
      RECT 5.948 0.932 6.038 1.15 ;
      RECT 5.994 0.887 6.107 0.943 ;
      RECT 6.038 0.849 6.069 0.978 ;
      RECT 6.254 0.427 6.344 0.924 ;
      RECT 6.069 0.834 6.344 0.924 ;
      RECT 5.923 0.427 6.344 0.517 ;
      RECT 5.923 0.205 6.013 0.517 ;
      RECT 4.691 0.96 5.15 1.05 ;
      RECT 4.662 0.907 4.691 1.036 ;
      RECT 2.86 0.755 3.15 1.035 ;
      RECT 4.662 0.96 5.192 1.029 ;
      RECT 4.616 0.87 4.662 0.998 ;
      RECT 4.616 0.96 5.23 0.989 ;
      RECT 5.112 0.941 5.856 0.97 ;
      RECT 4.616 0.941 4.729 0.998 ;
      RECT 4.57 0.824 4.616 0.952 ;
      RECT 5.15 0.901 5.856 0.97 ;
      RECT 4.524 0.778 4.57 0.906 ;
      RECT 5.192 0.88 5.856 0.97 ;
      RECT 5.766 0.741 5.856 0.97 ;
      RECT 4.486 0.824 4.616 0.864 ;
      RECT 2.86 0.755 4.524 0.845 ;
      RECT 5.766 0.741 5.902 0.779 ;
      RECT 3.938 0.395 4.028 0.845 ;
      RECT 5.812 0.696 5.923 0.746 ;
      RECT 5.812 0.696 5.961 0.716 ;
      RECT 5.923 0.607 6.118 0.697 ;
      RECT 5.856 0.651 6.118 0.697 ;
      RECT 5.902 0.617 5.923 0.746 ;
      RECT 3.533 0.395 4.46 0.485 ;
      RECT 2.807 0.395 3.443 0.485 ;
      RECT 3.353 0.17 3.443 0.485 ;
      RECT 4.808 0.265 5.351 0.355 ;
      RECT 4.797 0.221 4.808 0.35 ;
      RECT 4.751 0.193 4.797 0.321 ;
      RECT 4.713 0.246 4.846 0.279 ;
      RECT 3.353 0.17 4.751 0.26 ;
      RECT 4.919 0.575 5.059 0.87 ;
      RECT 4.118 0.575 5.059 0.665 ;
      RECT 4.562 0.38 4.705 0.665 ;
      RECT 2.155 1.14 3.797 1.23 ;
      RECT 3.707 0.935 3.797 1.23 ;
      RECT 3.707 0.935 4.184 1.025 ;
      RECT 2.163 0.96 2.77 1.05 ;
      RECT 2.68 0.575 2.77 1.05 ;
      RECT 1.81 0.88 1.95 1.018 ;
      RECT 1.06 0.88 2.254 0.97 ;
      RECT 1.06 0.548 1.15 0.97 ;
      RECT 2.68 0.575 3.828 0.665 ;
      RECT 1.106 0.503 1.196 0.586 ;
      RECT 1.106 0.503 1.234 0.544 ;
      RECT 1.196 0.435 1.966 0.525 ;
      RECT 1.15 0.458 1.966 0.525 ;
      RECT 2.45 0.7 2.59 0.87 ;
      RECT 1.285 0.7 2.59 0.79 ;
      RECT 2.065 0.2 2.155 0.79 ;
      RECT 2.065 0.2 3.263 0.29 ;
      RECT 1.755 1.14 2.065 1.23 ;
      RECT 1.713 1.081 1.755 1.209 ;
      RECT 0.775 1.095 0.97 1.185 ;
      RECT 0.88 0.36 0.97 1.185 ;
      RECT 1.675 1.14 2.065 1.169 ;
      RECT 0.88 1.06 1.713 1.15 ;
      RECT 0.775 1.121 1.793 1.15 ;
      RECT 0.88 0.36 1.02 0.45 ;
      RECT 0.045 0.915 0.185 1.11 ;
      RECT 0.045 0.915 0.79 1.005 ;
      RECT 0.7 0.795 0.79 1.005 ;
      RECT 0.045 0.25 0.135 1.11 ;
      RECT 0.045 0.283 0.727 0.373 ;
      RECT 0.637 0.17 0.727 0.373 ;
      RECT 0.045 0.25 0.185 0.373 ;
      RECT 0.637 0.17 1.172 0.26 ;
      RECT 0.7 0.473 0.79 0.635 ;
      RECT 0.226 0.473 0.366 0.585 ;
      RECT 0.226 0.473 0.79 0.563 ;
  END
END DFFSRQX1H7R

MACRO DFFSRQX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRQX2H7R 0 0 ;
  SIZE 7 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7 1.48 ;
        RECT 6.181 1.095 6.321 1.48 ;
        RECT 5.209 1.24 5.349 1.48 ;
        RECT 4.354 1.24 4.494 1.48 ;
        RECT 1.465 1.24 1.605 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7 0.08 ;
        RECT 6.181 -0.08 6.321 0.305 ;
        RECT 5.436 -0.08 5.576 0.175 ;
        RECT 1.455 -0.08 1.545 0.315 ;
        RECT 0.31 -0.08 0.45 0.193 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.66 0.25 1.975 0.345 ;
      LAYER MET2 ;
        RECT 1.85 0.18 1.95 0.56 ;
      LAYER VIA1 ;
        RECT 1.855 0.255 1.945 0.345 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.655 0.585 0.825 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.467 0.225 6.557 0.972 ;
        RECT 6.451 0.225 6.557 0.375 ;
      LAYER MET2 ;
        RECT 6.45 0.18 6.55 0.56 ;
      LAYER VIA1 ;
        RECT 6.455 0.255 6.545 0.345 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.015 0.567 5.145 0.776 ;
      LAYER MET2 ;
        RECT 5.05 0.43 5.15 0.96 ;
      LAYER VIA1 ;
        RECT 5.055 0.655 5.145 0.745 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.425 0.655 5.666 0.752 ;
        RECT 5.576 0.612 5.666 0.752 ;
      LAYER MET2 ;
        RECT 5.45 0.425 5.55 0.96 ;
      LAYER VIA1 ;
        RECT 5.455 0.655 5.545 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 4.614 1.14 5.091 1.23 ;
      RECT 3.887 1.14 4.235 1.23 ;
      RECT 4.572 1.14 5.133 1.209 ;
      RECT 3.887 1.14 4.277 1.209 ;
      RECT 5.931 1.06 6.071 1.18 ;
      RECT 5.981 0.834 6.071 1.18 ;
      RECT 4.534 1.14 5.171 1.169 ;
      RECT 3.887 1.14 4.315 1.169 ;
      RECT 5.133 1.06 6.071 1.15 ;
      RECT 5.053 1.121 6.071 1.15 ;
      RECT 5.091 1.081 5.133 1.209 ;
      RECT 4.197 1.121 4.652 1.15 ;
      RECT 4.235 1.081 4.614 1.15 ;
      RECT 4.277 1.06 4.572 1.15 ;
      RECT 5.981 0.834 6.377 0.924 ;
      RECT 6.287 0.427 6.377 0.924 ;
      RECT 5.956 0.427 6.377 0.517 ;
      RECT 5.956 0.205 6.046 0.517 ;
      RECT 4.691 0.96 5.015 1.05 ;
      RECT 4.662 0.907 4.691 1.036 ;
      RECT 2.86 0.755 3.35 1.035 ;
      RECT 4.662 0.96 5.057 1.029 ;
      RECT 4.616 0.87 4.662 0.998 ;
      RECT 4.616 0.96 5.095 0.989 ;
      RECT 5.797 0.607 5.887 0.97 ;
      RECT 4.977 0.941 5.887 0.97 ;
      RECT 5.057 0.88 5.887 0.97 ;
      RECT 4.616 0.941 4.729 0.998 ;
      RECT 4.57 0.824 4.616 0.952 ;
      RECT 5.015 0.901 5.887 0.97 ;
      RECT 4.524 0.778 4.57 0.906 ;
      RECT 4.486 0.824 4.616 0.864 ;
      RECT 2.86 0.755 4.524 0.845 ;
      RECT 3.938 0.395 4.028 0.845 ;
      RECT 5.797 0.607 6.151 0.697 ;
      RECT 3.543 0.395 4.46 0.485 ;
      RECT 2.807 0.395 3.453 0.485 ;
      RECT 3.363 0.215 3.453 0.485 ;
      RECT 5.701 0.295 5.841 0.47 ;
      RECT 5.39 0.295 5.841 0.385 ;
      RECT 5.349 0.236 5.39 0.365 ;
      RECT 5.303 0.193 5.349 0.321 ;
      RECT 3.363 0.215 4.632 0.305 ;
      RECT 5.303 0.276 5.428 0.321 ;
      RECT 5.265 0.17 5.303 0.279 ;
      RECT 4.546 0.17 5.303 0.26 ;
      RECT 4.784 0.38 4.924 0.87 ;
      RECT 4.118 0.575 4.924 0.665 ;
      RECT 4.784 0.38 5.257 0.47 ;
      RECT 2.155 1.14 3.797 1.23 ;
      RECT 3.707 0.935 3.797 1.23 ;
      RECT 3.707 0.935 4.184 1.025 ;
      RECT 2.163 0.96 2.77 1.05 ;
      RECT 2.68 0.575 2.77 1.05 ;
      RECT 1.81 0.88 1.95 1.018 ;
      RECT 1.06 0.88 2.254 0.97 ;
      RECT 1.06 0.548 1.15 0.97 ;
      RECT 2.68 0.575 3.848 0.665 ;
      RECT 1.106 0.503 1.196 0.586 ;
      RECT 1.106 0.503 1.234 0.544 ;
      RECT 1.196 0.435 1.966 0.525 ;
      RECT 1.15 0.458 1.966 0.525 ;
      RECT 2.45 0.7 2.59 0.87 ;
      RECT 1.285 0.7 2.59 0.79 ;
      RECT 2.065 0.2 2.155 0.79 ;
      RECT 2.065 0.2 3.273 0.29 ;
      RECT 1.755 1.14 2.065 1.23 ;
      RECT 1.713 1.081 1.755 1.209 ;
      RECT 0.775 1.095 0.97 1.185 ;
      RECT 0.88 0.36 0.97 1.185 ;
      RECT 1.675 1.14 2.065 1.169 ;
      RECT 0.88 1.06 1.713 1.15 ;
      RECT 0.775 1.121 1.793 1.15 ;
      RECT 0.88 0.36 1.02 0.45 ;
      RECT 0.045 0.915 0.185 1.11 ;
      RECT 0.045 0.915 0.79 1.005 ;
      RECT 0.7 0.795 0.79 1.005 ;
      RECT 0.045 0.25 0.135 1.11 ;
      RECT 0.045 0.283 0.727 0.373 ;
      RECT 0.637 0.17 0.727 0.373 ;
      RECT 0.045 0.25 0.185 0.373 ;
      RECT 0.637 0.17 1.172 0.26 ;
      RECT 0.7 0.473 0.79 0.635 ;
      RECT 0.226 0.473 0.366 0.585 ;
      RECT 0.226 0.473 0.79 0.563 ;
  END
END DFFSRQX2H7R

MACRO DFFSRX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRX0P5H7R 0 0 ;
  SIZE 6.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.2 1.48 ;
        RECT 5.715 1.24 5.855 1.48 ;
        RECT 5.195 1.24 5.335 1.48 ;
        RECT 4.385 1.24 4.525 1.48 ;
        RECT 3.76 1.24 3.9 1.48 ;
        RECT 1.345 1.235 1.485 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.2 0.08 ;
        RECT 5.765 -0.08 5.855 0.33 ;
        RECT 5.28 -0.08 5.37 0.33 ;
        RECT 4.505 -0.08 4.645 0.16 ;
        RECT 1.38 -0.08 1.52 0.16 ;
        RECT 0.36 -0.08 0.5 0.16 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.865 0.75 2.145 0.84 ;
        RECT 2.055 0.625 2.145 0.84 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.655 0.575 0.82 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.015 0.425 6.145 0.575 ;
        RECT 6.015 0.245 6.105 1.045 ;
      LAYER MET2 ;
        RECT 6.05 0.23 6.15 0.76 ;
      LAYER VIA1 ;
        RECT 6.055 0.455 6.145 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.455 0.88 5.65 0.97 ;
        RECT 5.535 0.255 5.625 0.6 ;
        RECT 5.455 0.51 5.545 0.97 ;
      LAYER MET2 ;
        RECT 5.45 0.425 5.55 0.96 ;
      LAYER VIA1 ;
        RECT 5.455 0.655 5.545 0.745 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.395 0.455 4.575 0.545 ;
        RECT 4.355 0.52 4.51 0.61 ;
      LAYER MET2 ;
        RECT 4.45 0.225 4.55 0.76 ;
      LAYER VIA1 ;
        RECT 4.455 0.455 4.545 0.545 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.585 0.67 4.775 0.785 ;
        RECT 4.655 0.625 4.775 0.785 ;
      LAYER MET2 ;
        RECT 4.65 0.425 4.75 0.96 ;
      LAYER VIA1 ;
        RECT 4.655 0.655 4.745 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 3.225 1.14 3.607 1.23 ;
      RECT 4.88 1.06 5.02 1.185 ;
      RECT 5.74 0.615 5.83 1.15 ;
      RECT 3.517 1.06 5.83 1.15 ;
      RECT 5.1 0.295 5.19 1.15 ;
      RECT 5 0.295 5.19 0.385 ;
      RECT 2.845 0.873 2.935 1.05 ;
      RECT 4.345 0.88 5.01 0.97 ;
      RECT 4.92 0.56 5.01 0.97 ;
      RECT 4.345 0.7 4.435 0.97 ;
      RECT 2.891 0.828 2.981 0.911 ;
      RECT 2.891 0.828 3.019 0.869 ;
      RECT 3.415 0.439 3.505 0.85 ;
      RECT 2.935 0.783 3.505 0.85 ;
      RECT 2.981 0.76 3.505 0.85 ;
      RECT 3.415 0.7 4.435 0.79 ;
      RECT 3.415 0.475 3.799 0.565 ;
      RECT 3.415 0.475 3.856 0.531 ;
      RECT 3.394 0.36 3.415 0.489 ;
      RECT 3.81 0.35 3.902 0.485 ;
      RECT 3.761 0.456 3.902 0.485 ;
      RECT 3.799 0.431 3.81 0.56 ;
      RECT 3.356 0.439 3.505 0.459 ;
      RECT 3.799 0.431 3.924 0.451 ;
      RECT 3.81 0.35 3.95 0.44 ;
      RECT 3.07 0.35 3.394 0.44 ;
      RECT 3.07 0.394 3.461 0.44 ;
      RECT 3.545 0.17 3.685 0.36 ;
      RECT 4.436 0.26 4.885 0.35 ;
      RECT 4.795 0.21 4.885 0.35 ;
      RECT 4.43 0.219 4.436 0.347 ;
      RECT 4.384 0.193 4.43 0.321 ;
      RECT 4.346 0.26 4.885 0.279 ;
      RECT 2.42 0.17 4.384 0.26 ;
      RECT 2.42 0.241 4.474 0.26 ;
      RECT 3.995 0.52 4.145 0.61 ;
      RECT 4.055 0.35 4.145 0.61 ;
      RECT 4.055 0.35 4.305 0.44 ;
      RECT 1.98 1.14 3.135 1.23 ;
      RECT 3.045 0.993 3.135 1.23 ;
      RECT 3.091 0.955 3.135 1.23 ;
      RECT 1.98 1.125 2.12 1.23 ;
      RECT 3.045 0.993 3.159 1.042 ;
      RECT 3.121 0.94 3.42 1.03 ;
      RECT 2.209 0.96 2.58 1.05 ;
      RECT 2.49 0.825 2.58 1.05 ;
      RECT 2.171 0.935 2.184 1.05 ;
      RECT 1.694 0.935 2.146 1.025 ;
      RECT 1.025 0.835 1.095 0.995 ;
      RECT 1.185 0.875 1.616 0.965 ;
      RECT 1.694 0.915 1.8 1.025 ;
      RECT 2.49 0.825 2.641 0.915 ;
      RECT 2.954 0.55 3.325 0.64 ;
      RECT 1.234 0.43 1.635 0.52 ;
      RECT 1.733 0.37 1.835 0.46 ;
      RECT 2.916 0.55 2.954 0.659 ;
      RECT 2.909 0.553 2.916 0.682 ;
      RECT 2.863 0.58 2.909 0.708 ;
      RECT 2.817 0.626 2.863 0.754 ;
      RECT 2.771 0.672 2.817 0.8 ;
      RECT 2.725 0.718 2.771 0.846 ;
      RECT 2.679 0.764 2.725 0.892 ;
      RECT 2.641 0.806 2.679 0.915 ;
      RECT 2.184 0.947 2.209 1.05 ;
      RECT 2.146 0.935 2.171 1.038 ;
      RECT 1.695 0.37 1.733 0.479 ;
      RECT 1.673 0.381 1.695 0.509 ;
      RECT 1.676 0.906 1.694 1.025 ;
      RECT 1.654 0.886 1.676 1.014 ;
      RECT 1.635 0.411 1.673 0.52 ;
      RECT 1.616 0.875 1.654 0.984 ;
      RECT 1.196 0.43 1.234 0.539 ;
      RECT 1.185 0.435 1.196 0.564 ;
      RECT 1.161 0.453 1.185 0.965 ;
      RECT 1.115 0.488 1.161 0.965 ;
      RECT 1.095 0.521 1.115 0.995 ;
      RECT 2.26 0.78 2.4 0.87 ;
      RECT 2.26 0.563 2.35 0.87 ;
      RECT 1.275 0.61 1.756 0.7 ;
      RECT 1.275 0.61 1.771 0.693 ;
      RECT 1.275 0.61 1.809 0.666 ;
      RECT 2.26 0.563 2.676 0.653 ;
      RECT 1.275 0.61 1.904 0.647 ;
      RECT 2.26 0.563 2.722 0.63 ;
      RECT 1.718 0.591 1.95 0.624 ;
      RECT 2.221 0.464 2.26 0.593 ;
      RECT 1.756 0.564 1.955 0.599 ;
      RECT 1.771 0.557 2.001 0.573 ;
      RECT 1.95 0.47 1.955 0.599 ;
      RECT 2.638 0.544 2.781 0.571 ;
      RECT 2.722 0.472 2.735 0.601 ;
      RECT 2.221 0.546 2.339 0.593 ;
      RECT 1.866 0.538 2.001 0.573 ;
      RECT 1.904 0.496 1.95 0.624 ;
      RECT 2.183 0.507 2.306 0.554 ;
      RECT 2.676 0.502 2.781 0.571 ;
      RECT 1.955 0.35 2.016 0.543 ;
      RECT 1.955 0.445 2.221 0.535 ;
      RECT 2.735 0.35 2.825 0.526 ;
      RECT 1.955 0.35 2.045 0.535 ;
      RECT 0.045 0.915 0.185 1.025 ;
      RECT 0.045 0.915 0.755 1.005 ;
      RECT 0.665 0.74 0.755 1.005 ;
      RECT 0.045 0.265 0.135 1.025 ;
      RECT 2.369 0.375 2.594 0.465 ;
      RECT 2.33 0.317 2.369 0.446 ;
      RECT 2.286 0.356 2.407 0.404 ;
      RECT 2.24 0.17 2.33 0.359 ;
      RECT 0.045 0.265 0.685 0.355 ;
      RECT 0.595 0.17 0.685 0.355 ;
      RECT 1.19 0.25 1.596 0.34 ;
      RECT 1.19 0.25 1.676 0.279 ;
      RECT 1.638 0.17 2.33 0.26 ;
      RECT 1.558 0.231 2.33 0.26 ;
      RECT 1.596 0.191 1.638 0.319 ;
      RECT 0.595 0.17 1.28 0.26 ;
      RECT 1.62 1.14 1.89 1.23 ;
      RECT 1.574 1.078 1.62 1.206 ;
      RECT 0.755 1.095 1.229 1.185 ;
      RECT 1.536 1.14 1.89 1.164 ;
      RECT 0.755 1.095 1.269 1.164 ;
      RECT 1.231 1.055 1.574 1.145 ;
      RECT 0.755 1.121 1.659 1.145 ;
      RECT 0.755 1.101 1.621 1.145 ;
      RECT 1.229 1.056 1.231 1.184 ;
      RECT 0.845 0.733 0.935 1.185 ;
      RECT 1.191 1.076 1.574 1.145 ;
      RECT 0.845 0.733 0.981 0.771 ;
      RECT 0.915 0.363 1.005 0.736 ;
      RECT 0.891 0.698 1.005 0.736 ;
      RECT 0.89 0.363 1.03 0.453 ;
      RECT 0.73 0.492 0.82 0.65 ;
      RECT 0.225 0.475 0.315 0.645 ;
      RECT 0.225 0.475 0.785 0.565 ;
      RECT 3.865 0.88 4.21 0.97 ;
  END
END DFFSRX0P5H7R

MACRO DFFSRX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRX1H7R 0 0 ;
  SIZE 6.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.2 1.48 ;
        RECT 5.715 1.24 5.855 1.48 ;
        RECT 5.195 1.24 5.335 1.48 ;
        RECT 4.385 1.24 4.525 1.48 ;
        RECT 3.76 1.24 3.9 1.48 ;
        RECT 1.345 1.235 1.485 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.2 0.08 ;
        RECT 5.765 -0.08 5.855 0.33 ;
        RECT 5.28 -0.08 5.37 0.33 ;
        RECT 4.505 -0.08 4.645 0.16 ;
        RECT 1.38 -0.08 1.52 0.16 ;
        RECT 0.36 -0.08 0.5 0.16 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.865 0.75 2.145 0.84 ;
        RECT 2.055 0.625 2.145 0.84 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.655 0.575 0.82 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.015 0.295 6.145 1.19 ;
      LAYER MET2 ;
        RECT 6.05 0.23 6.15 0.76 ;
      LAYER VIA1 ;
        RECT 6.055 0.455 6.145 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.455 0.825 5.65 0.915 ;
        RECT 5.535 0.265 5.625 0.6 ;
        RECT 5.455 0.51 5.545 0.915 ;
      LAYER MET2 ;
        RECT 5.45 0.425 5.55 0.96 ;
      LAYER VIA1 ;
        RECT 5.455 0.655 5.545 0.745 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.395 0.455 4.575 0.545 ;
        RECT 4.355 0.52 4.51 0.61 ;
      LAYER MET2 ;
        RECT 4.45 0.225 4.55 0.76 ;
      LAYER VIA1 ;
        RECT 4.455 0.455 4.545 0.545 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.585 0.67 4.775 0.785 ;
        RECT 4.655 0.625 4.775 0.785 ;
      LAYER MET2 ;
        RECT 4.65 0.425 4.75 0.96 ;
      LAYER VIA1 ;
        RECT 4.655 0.655 4.745 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 3.225 1.14 3.607 1.23 ;
      RECT 4.88 1.06 5.02 1.185 ;
      RECT 3.517 1.06 5.674 1.15 ;
      RECT 3.517 1.06 5.72 1.127 ;
      RECT 5.636 1.041 5.786 1.061 ;
      RECT 5.72 0.966 5.74 1.094 ;
      RECT 5.1 0.3 5.19 1.15 ;
      RECT 5.674 0.999 5.786 1.061 ;
      RECT 5.74 0.615 5.83 1.016 ;
      RECT 5 0.3 5.19 0.39 ;
      RECT 2.845 0.873 2.935 1.05 ;
      RECT 4.345 0.88 5.01 0.97 ;
      RECT 4.92 0.56 5.01 0.97 ;
      RECT 4.345 0.7 4.435 0.97 ;
      RECT 2.891 0.828 2.981 0.911 ;
      RECT 2.891 0.828 3.019 0.869 ;
      RECT 3.415 0.43 3.505 0.85 ;
      RECT 2.935 0.783 3.505 0.85 ;
      RECT 2.981 0.76 3.505 0.85 ;
      RECT 3.415 0.7 4.435 0.79 ;
      RECT 3.415 0.43 3.764 0.52 ;
      RECT 3.415 0.43 3.844 0.459 ;
      RECT 3.381 0.43 3.844 0.457 ;
      RECT 3.806 0.35 3.95 0.44 ;
      RECT 3.726 0.411 3.95 0.44 ;
      RECT 3.764 0.371 3.806 0.499 ;
      RECT 3.07 0.413 3.499 0.44 ;
      RECT 3.07 0.373 3.465 0.44 ;
      RECT 3.07 0.35 3.419 0.44 ;
      RECT 4.436 0.26 4.885 0.35 ;
      RECT 4.795 0.21 4.885 0.35 ;
      RECT 4.43 0.219 4.436 0.347 ;
      RECT 3.545 0.17 3.685 0.34 ;
      RECT 4.384 0.193 4.43 0.321 ;
      RECT 4.346 0.26 4.885 0.279 ;
      RECT 2.42 0.17 4.384 0.26 ;
      RECT 2.42 0.241 4.474 0.26 ;
      RECT 3.995 0.52 4.145 0.61 ;
      RECT 4.055 0.35 4.145 0.61 ;
      RECT 4.055 0.35 4.305 0.44 ;
      RECT 1.98 1.14 3.135 1.23 ;
      RECT 3.045 0.993 3.135 1.23 ;
      RECT 3.091 0.955 3.135 1.23 ;
      RECT 1.98 1.125 2.12 1.23 ;
      RECT 3.045 0.993 3.159 1.042 ;
      RECT 3.121 0.94 3.42 1.03 ;
      RECT 2.209 0.96 2.58 1.05 ;
      RECT 2.49 0.825 2.58 1.05 ;
      RECT 2.171 0.935 2.184 1.05 ;
      RECT 1.694 0.935 2.146 1.025 ;
      RECT 1.025 0.835 1.095 0.995 ;
      RECT 1.185 0.875 1.616 0.965 ;
      RECT 1.694 0.915 1.8 1.025 ;
      RECT 2.49 0.825 2.641 0.915 ;
      RECT 2.954 0.55 3.325 0.64 ;
      RECT 1.234 0.43 1.635 0.52 ;
      RECT 1.733 0.37 1.835 0.46 ;
      RECT 2.916 0.55 2.954 0.659 ;
      RECT 2.909 0.553 2.916 0.682 ;
      RECT 2.863 0.58 2.909 0.708 ;
      RECT 2.817 0.626 2.863 0.754 ;
      RECT 2.771 0.672 2.817 0.8 ;
      RECT 2.725 0.718 2.771 0.846 ;
      RECT 2.679 0.764 2.725 0.892 ;
      RECT 2.641 0.806 2.679 0.915 ;
      RECT 2.184 0.947 2.209 1.05 ;
      RECT 2.146 0.935 2.171 1.038 ;
      RECT 1.695 0.37 1.733 0.479 ;
      RECT 1.673 0.381 1.695 0.509 ;
      RECT 1.676 0.906 1.694 1.025 ;
      RECT 1.654 0.886 1.676 1.014 ;
      RECT 1.635 0.411 1.673 0.52 ;
      RECT 1.616 0.875 1.654 0.984 ;
      RECT 1.196 0.43 1.234 0.539 ;
      RECT 1.185 0.435 1.196 0.564 ;
      RECT 1.161 0.453 1.185 0.965 ;
      RECT 1.115 0.488 1.161 0.965 ;
      RECT 1.095 0.521 1.115 0.995 ;
      RECT 2.26 0.78 2.4 0.87 ;
      RECT 2.26 0.563 2.35 0.87 ;
      RECT 1.275 0.61 1.756 0.7 ;
      RECT 1.275 0.61 1.771 0.693 ;
      RECT 1.275 0.61 1.809 0.666 ;
      RECT 2.26 0.563 2.676 0.653 ;
      RECT 1.275 0.61 1.904 0.647 ;
      RECT 2.26 0.563 2.722 0.63 ;
      RECT 1.718 0.591 1.95 0.624 ;
      RECT 2.221 0.464 2.26 0.593 ;
      RECT 1.756 0.564 1.955 0.599 ;
      RECT 1.771 0.557 2.001 0.573 ;
      RECT 1.95 0.47 1.955 0.599 ;
      RECT 2.638 0.544 2.781 0.571 ;
      RECT 2.722 0.472 2.735 0.601 ;
      RECT 2.221 0.546 2.339 0.593 ;
      RECT 1.866 0.538 2.001 0.573 ;
      RECT 1.904 0.496 1.95 0.624 ;
      RECT 2.183 0.507 2.306 0.554 ;
      RECT 2.676 0.502 2.781 0.571 ;
      RECT 1.955 0.35 2.016 0.543 ;
      RECT 1.955 0.445 2.221 0.535 ;
      RECT 2.735 0.35 2.825 0.526 ;
      RECT 1.955 0.35 2.045 0.535 ;
      RECT 0.045 0.915 0.185 1.025 ;
      RECT 0.045 0.915 0.755 1.005 ;
      RECT 0.665 0.74 0.755 1.005 ;
      RECT 0.045 0.265 0.135 1.025 ;
      RECT 2.369 0.375 2.594 0.465 ;
      RECT 2.33 0.317 2.369 0.446 ;
      RECT 2.286 0.356 2.407 0.404 ;
      RECT 2.24 0.17 2.33 0.359 ;
      RECT 0.045 0.265 0.685 0.355 ;
      RECT 0.595 0.17 0.685 0.355 ;
      RECT 1.19 0.25 1.596 0.34 ;
      RECT 1.19 0.25 1.676 0.279 ;
      RECT 1.638 0.17 2.33 0.26 ;
      RECT 1.558 0.231 2.33 0.26 ;
      RECT 1.596 0.191 1.638 0.319 ;
      RECT 0.595 0.17 1.28 0.26 ;
      RECT 1.62 1.14 1.89 1.23 ;
      RECT 1.574 1.078 1.62 1.206 ;
      RECT 0.755 1.095 1.229 1.185 ;
      RECT 1.536 1.14 1.89 1.164 ;
      RECT 0.755 1.095 1.269 1.164 ;
      RECT 1.231 1.055 1.574 1.145 ;
      RECT 0.755 1.121 1.659 1.145 ;
      RECT 0.755 1.101 1.621 1.145 ;
      RECT 1.229 1.056 1.231 1.184 ;
      RECT 0.845 0.733 0.935 1.185 ;
      RECT 1.191 1.076 1.574 1.145 ;
      RECT 0.845 0.733 0.981 0.771 ;
      RECT 0.915 0.363 1.005 0.736 ;
      RECT 0.891 0.698 1.005 0.736 ;
      RECT 0.89 0.363 1.03 0.453 ;
      RECT 0.73 0.492 0.82 0.65 ;
      RECT 0.225 0.475 0.315 0.645 ;
      RECT 0.225 0.475 0.785 0.565 ;
      RECT 3.865 0.88 4.21 0.97 ;
  END
END DFFSRX1H7R

MACRO DFFSRX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRX2H7R 0 0 ;
  SIZE 6.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.4 1.48 ;
        RECT 5.69 1.215 5.78 1.48 ;
        RECT 5.145 1.24 5.285 1.48 ;
        RECT 4.335 1.24 4.475 1.48 ;
        RECT 3.715 1.24 3.855 1.48 ;
        RECT 1.345 1.235 1.485 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.4 0.08 ;
        RECT 5.715 -0.08 5.805 0.33 ;
        RECT 5.235 -0.08 5.325 0.33 ;
        RECT 4.46 -0.08 4.6 0.16 ;
        RECT 1.38 -0.08 1.52 0.16 ;
        RECT 0.36 -0.08 0.5 0.16 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.865 0.75 2.145 0.84 ;
        RECT 2.055 0.625 2.145 0.84 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.655 0.575 0.82 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.005 0.805 6.145 1.145 ;
        RECT 6.055 0.36 6.145 1.145 ;
        RECT 5.945 0.36 6.145 0.45 ;
      LAYER MET2 ;
        RECT 6.05 0.23 6.15 0.76 ;
      LAYER VIA1 ;
        RECT 6.055 0.455 6.145 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.455 0.36 5.61 0.45 ;
        RECT 5.455 0.825 5.6 0.915 ;
        RECT 5.455 0.36 5.545 0.915 ;
      LAYER MET2 ;
        RECT 5.45 0.225 5.55 0.76 ;
      LAYER VIA1 ;
        RECT 5.455 0.455 5.545 0.545 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.35 0.455 4.575 0.545 ;
        RECT 4.305 0.52 4.45 0.61 ;
      LAYER MET2 ;
        RECT 4.45 0.225 4.55 0.76 ;
      LAYER VIA1 ;
        RECT 4.455 0.455 4.545 0.545 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.535 0.67 4.745 0.785 ;
        RECT 4.655 0.625 4.745 0.785 ;
      LAYER MET2 ;
        RECT 4.65 0.425 4.75 0.96 ;
      LAYER VIA1 ;
        RECT 4.655 0.655 4.745 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 3.135 1.14 3.562 1.23 ;
      RECT 4.83 1.06 4.97 1.185 ;
      RECT 3.472 1.06 5.624 1.15 ;
      RECT 3.472 1.06 5.67 1.127 ;
      RECT 5.586 1.041 5.736 1.061 ;
      RECT 5.67 0.966 5.69 1.094 ;
      RECT 5.05 0.32 5.14 1.15 ;
      RECT 5.624 0.999 5.736 1.061 ;
      RECT 5.69 0.615 5.78 1.016 ;
      RECT 4.96 0.32 5.14 0.41 ;
      RECT 2.775 0.76 2.865 1.05 ;
      RECT 4.295 0.88 4.96 0.97 ;
      RECT 4.87 0.56 4.96 0.97 ;
      RECT 4.295 0.7 4.385 0.97 ;
      RECT 2.775 0.76 3.46 0.85 ;
      RECT 3.37 0.41 3.46 0.85 ;
      RECT 3.37 0.7 4.385 0.79 ;
      RECT 3.37 0.41 3.739 0.5 ;
      RECT 3.37 0.41 3.799 0.459 ;
      RECT 3.336 0.41 3.799 0.457 ;
      RECT 3.761 0.35 3.905 0.44 ;
      RECT 3.701 0.391 3.905 0.44 ;
      RECT 3.739 0.361 3.761 0.489 ;
      RECT 3.025 0.403 3.434 0.44 ;
      RECT 3.025 0.373 3.42 0.44 ;
      RECT 3.025 0.35 3.374 0.44 ;
      RECT 4.391 0.26 4.84 0.35 ;
      RECT 4.75 0.21 4.84 0.35 ;
      RECT 4.385 0.219 4.391 0.347 ;
      RECT 4.339 0.193 4.385 0.321 ;
      RECT 3.5 0.17 3.64 0.32 ;
      RECT 2.185 0.17 2.325 0.29 ;
      RECT 4.301 0.26 4.84 0.279 ;
      RECT 2.185 0.17 4.339 0.26 ;
      RECT 2.185 0.241 4.429 0.26 ;
      RECT 3.95 0.52 4.095 0.61 ;
      RECT 4.005 0.35 4.095 0.61 ;
      RECT 4.005 0.35 4.26 0.44 ;
      RECT 1.98 1.14 3.045 1.23 ;
      RECT 2.955 0.94 3.045 1.23 ;
      RECT 1.98 1.115 2.12 1.23 ;
      RECT 2.955 0.94 3.375 1.03 ;
      RECT 2.776 0.55 3.28 0.64 ;
      RECT 2.751 0.55 3.28 0.628 ;
      RECT 2.705 0.425 2.795 0.592 ;
      RECT 2.705 0.54 2.814 0.592 ;
      RECT 2.45 0.96 2.685 1.05 ;
      RECT 2.595 0.669 2.685 1.05 ;
      RECT 2.571 0.669 2.685 0.707 ;
      RECT 1.275 0.61 1.761 0.7 ;
      RECT 1.275 0.61 1.776 0.693 ;
      RECT 2.525 0.415 2.615 0.672 ;
      RECT 2.525 0.634 2.661 0.672 ;
      RECT 1.275 0.61 1.814 0.666 ;
      RECT 1.275 0.61 1.904 0.647 ;
      RECT 1.723 0.591 1.92 0.639 ;
      RECT 1.761 0.564 1.966 0.608 ;
      RECT 1.904 0.511 1.92 0.639 ;
      RECT 1.776 0.557 1.966 0.608 ;
      RECT 1.866 0.538 1.904 0.647 ;
      RECT 1.92 0.415 2.01 0.563 ;
      RECT 1.92 0.415 2.615 0.505 ;
      RECT 1.746 0.935 2.335 1.025 ;
      RECT 2.245 0.76 2.335 1.025 ;
      RECT 1.732 0.935 2.335 1.018 ;
      RECT 1.025 0.835 1.115 0.995 ;
      RECT 1.686 0.935 2.335 0.988 ;
      RECT 1.025 0.875 1.77 0.965 ;
      RECT 1.025 0.928 1.784 0.965 ;
      RECT 2.245 0.76 2.505 0.85 ;
      RECT 1.095 0.521 1.185 0.965 ;
      RECT 1.115 0.488 1.234 0.539 ;
      RECT 1.185 0.435 1.196 0.564 ;
      RECT 1.115 0.488 1.673 0.52 ;
      RECT 1.161 0.453 1.69 0.512 ;
      RECT 1.161 0.453 1.728 0.484 ;
      RECT 1.69 0.375 1.83 0.465 ;
      RECT 1.673 0.383 1.69 0.512 ;
      RECT 1.196 0.43 1.83 0.465 ;
      RECT 1.635 0.411 1.673 0.52 ;
      RECT 0.045 0.915 0.755 1.005 ;
      RECT 0.665 0.74 0.755 1.005 ;
      RECT 0.045 0.265 0.135 1.005 ;
      RECT 0.045 0.265 0.685 0.355 ;
      RECT 0.595 0.17 0.685 0.355 ;
      RECT 1.19 0.25 1.596 0.34 ;
      RECT 1.19 0.25 1.676 0.279 ;
      RECT 1.638 0.17 1.915 0.26 ;
      RECT 1.558 0.231 1.915 0.26 ;
      RECT 1.596 0.191 1.638 0.319 ;
      RECT 0.595 0.17 1.28 0.26 ;
      RECT 1.62 1.14 1.89 1.23 ;
      RECT 1.574 1.078 1.62 1.206 ;
      RECT 0.755 1.095 1.229 1.185 ;
      RECT 1.536 1.14 1.89 1.164 ;
      RECT 0.755 1.095 1.269 1.164 ;
      RECT 1.231 1.055 1.574 1.145 ;
      RECT 0.755 1.121 1.659 1.145 ;
      RECT 0.755 1.101 1.621 1.145 ;
      RECT 1.229 1.056 1.231 1.184 ;
      RECT 0.845 0.733 0.935 1.185 ;
      RECT 1.191 1.076 1.574 1.145 ;
      RECT 0.845 0.733 0.981 0.771 ;
      RECT 0.915 0.363 1.005 0.736 ;
      RECT 0.891 0.698 1.005 0.736 ;
      RECT 0.89 0.363 1.03 0.453 ;
      RECT 0.73 0.492 0.82 0.65 ;
      RECT 0.225 0.475 0.315 0.645 ;
      RECT 0.225 0.475 0.785 0.565 ;
      RECT 3.82 0.88 4.16 0.97 ;
  END
END DFFSRX2H7R

MACRO DFFSX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSX0P5H7R 0 0 ;
  SIZE 5.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.6 1.48 ;
        RECT 5.317 1.055 5.407 1.48 ;
        RECT 4.387 1.225 4.527 1.48 ;
        RECT 3.555 1.225 3.695 1.48 ;
        RECT 2.312 1.225 2.452 1.48 ;
        RECT 1.46 1.225 1.6 1.48 ;
        RECT 0.31 1.14 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.6 0.08 ;
        RECT 4.807 -0.08 4.897 0.347 ;
        RECT 4.307 -0.08 4.397 0.33 ;
        RECT 3.802 -0.08 3.942 0.34 ;
        RECT 1.42 -0.08 1.56 0.175 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.425 0.345 0.65 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.6 0.545 0.87 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.067 0.225 5.157 1.066 ;
        RECT 5.035 0.225 5.157 0.375 ;
      LAYER MET2 ;
        RECT 5.05 0.18 5.15 0.56 ;
      LAYER VIA1 ;
        RECT 5.055 0.255 5.145 0.345 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.625 0.855 4.792 0.945 ;
        RECT 4.625 0.28 4.715 0.945 ;
        RECT 4.527 0.28 4.715 0.37 ;
      LAYER MET2 ;
        RECT 4.65 0.625 4.75 1.16 ;
      LAYER VIA1 ;
        RECT 4.655 0.855 4.745 0.945 ;
    END
  END QN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.65 0.625 3.785 0.825 ;
      LAYER MET2 ;
        RECT 3.65 0.43 3.75 0.96 ;
      LAYER VIA1 ;
        RECT 3.655 0.655 3.745 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 3.462 1.045 4.977 1.135 ;
      RECT 4.887 0.551 4.977 1.135 ;
      RECT 4.445 0.468 4.535 1.135 ;
      RECT 3.462 0.655 3.552 1.135 ;
      RECT 4.108 0.468 4.535 0.558 ;
      RECT 4.103 0.468 4.535 0.556 ;
      RECT 4.057 0.255 4.147 0.53 ;
      RECT 2.877 0.89 3.038 0.98 ;
      RECT 2.948 0.355 3.038 0.98 ;
      RECT 3.907 0.557 3.997 0.955 ;
      RECT 3.907 0.648 4.355 0.738 ;
      RECT 3.907 0.636 4.066 0.738 ;
      RECT 3.907 0.602 4.043 0.738 ;
      RECT 3.894 0.482 3.907 0.611 ;
      RECT 3.848 0.453 3.894 0.581 ;
      RECT 3.848 0.512 3.953 0.581 ;
      RECT 3.81 0.512 3.953 0.539 ;
      RECT 2.948 0.43 3.848 0.52 ;
      RECT 2.948 0.355 3.088 0.52 ;
      RECT 3.552 0.17 3.692 0.34 ;
      RECT 2.1 0.17 3.692 0.26 ;
      RECT 2.585 1.14 3.347 1.23 ;
      RECT 1.733 1.14 2.148 1.23 ;
      RECT 0.69 1.14 1.199 1.23 ;
      RECT 2.574 1.096 2.585 1.225 ;
      RECT 1.722 1.096 1.733 1.225 ;
      RECT 2.528 1.068 2.574 1.196 ;
      RECT 1.676 1.068 1.722 1.196 ;
      RECT 3.232 0.655 3.322 1.23 ;
      RECT 2.49 1.121 2.623 1.154 ;
      RECT 2.11 1.121 2.243 1.154 ;
      RECT 2.194 1.05 2.205 1.179 ;
      RECT 1.638 1.121 1.771 1.154 ;
      RECT 1.161 1.121 1.294 1.154 ;
      RECT 1.245 1.05 1.256 1.179 ;
      RECT 0.69 0.465 0.78 1.23 ;
      RECT 2.205 1.045 2.528 1.135 ;
      RECT 1.256 1.045 1.676 1.135 ;
      RECT 2.148 1.079 2.194 1.207 ;
      RECT 1.199 1.079 1.245 1.207 ;
      RECT 0.045 0.96 0.78 1.05 ;
      RECT 0.045 0.252 0.135 1.05 ;
      RECT 0.045 0.252 0.185 0.342 ;
      RECT 2.652 0.71 2.742 0.991 ;
      RECT 2.652 0.71 2.858 0.8 ;
      RECT 2.768 0.35 2.858 0.8 ;
      RECT 1.255 0.505 2.037 0.595 ;
      RECT 1.947 0.35 2.037 0.595 ;
      RECT 1.947 0.35 2.858 0.44 ;
      RECT 1.87 0.685 2.01 0.855 ;
      RECT 1.05 0.685 2.22 0.775 ;
      RECT 2.13 0.53 2.22 0.775 ;
      RECT 1.05 0.325 1.14 0.775 ;
      RECT 2.13 0.53 2.678 0.62 ;
      RECT 1.05 0.325 1.857 0.415 ;
      RECT 1.767 0.205 1.857 0.415 ;
      RECT 1.809 0.96 2.071 1.05 ;
      RECT 1.798 0.916 1.809 1.045 ;
      RECT 0.87 0.245 0.96 1.03 ;
      RECT 1.798 0.96 2.117 1.027 ;
      RECT 1.752 0.888 1.798 1.016 ;
      RECT 2.033 0.941 2.166 0.974 ;
      RECT 2.117 0.87 2.128 0.999 ;
      RECT 1.714 0.941 1.847 0.974 ;
      RECT 2.128 0.865 2.33 0.955 ;
      RECT 0.87 0.865 1.752 0.955 ;
      RECT 2.071 0.899 2.33 0.955 ;
      RECT 0.805 0.245 0.96 0.335 ;
  END
END DFFSX0P5H7R

MACRO DFFSX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSX1H7R 0 0 ;
  SIZE 5.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.6 1.48 ;
        RECT 5.317 0.87 5.407 1.48 ;
        RECT 4.387 1.225 4.527 1.48 ;
        RECT 3.555 1.225 3.695 1.48 ;
        RECT 2.312 1.225 2.452 1.48 ;
        RECT 1.46 1.225 1.6 1.48 ;
        RECT 0.31 1.14 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.6 0.08 ;
        RECT 4.807 -0.08 4.897 0.347 ;
        RECT 4.307 -0.08 4.397 0.33 ;
        RECT 3.802 -0.08 3.942 0.34 ;
        RECT 1.42 -0.08 1.56 0.175 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.425 0.345 0.65 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.6 0.545 0.87 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.067 0.225 5.157 1.191 ;
        RECT 5.035 0.225 5.157 0.375 ;
      LAYER MET2 ;
        RECT 5.05 0.18 5.15 0.56 ;
      LAYER VIA1 ;
        RECT 5.055 0.255 5.145 0.345 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.625 0.855 4.792 0.945 ;
        RECT 4.625 0.232 4.715 0.945 ;
        RECT 4.527 0.232 4.715 0.322 ;
      LAYER MET2 ;
        RECT 4.65 0.625 4.75 1.16 ;
      LAYER VIA1 ;
        RECT 4.655 0.855 4.745 0.945 ;
    END
  END QN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.65 0.625 3.785 0.825 ;
      LAYER MET2 ;
        RECT 3.65 0.43 3.75 0.96 ;
      LAYER VIA1 ;
        RECT 3.655 0.655 3.745 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 3.462 1.045 4.977 1.135 ;
      RECT 4.887 0.551 4.977 1.135 ;
      RECT 4.445 0.42 4.535 1.135 ;
      RECT 3.462 0.655 3.552 1.135 ;
      RECT 4.105 0.42 4.535 0.51 ;
      RECT 4.103 0.42 4.535 0.509 ;
      RECT 4.057 0.275 4.147 0.485 ;
      RECT 2.877 0.89 3.038 0.98 ;
      RECT 2.948 0.355 3.038 0.98 ;
      RECT 3.907 0.557 3.997 0.955 ;
      RECT 3.907 0.6 4.355 0.69 ;
      RECT 3.894 0.482 3.907 0.611 ;
      RECT 3.894 0.589 4.018 0.611 ;
      RECT 3.848 0.453 3.894 0.581 ;
      RECT 3.848 0.512 3.953 0.581 ;
      RECT 3.81 0.512 3.953 0.539 ;
      RECT 2.948 0.43 3.848 0.52 ;
      RECT 2.948 0.355 3.088 0.52 ;
      RECT 3.552 0.17 3.692 0.34 ;
      RECT 2.1 0.17 3.692 0.26 ;
      RECT 2.585 1.14 3.347 1.23 ;
      RECT 1.733 1.14 2.148 1.23 ;
      RECT 0.69 1.14 1.199 1.23 ;
      RECT 2.574 1.096 2.585 1.225 ;
      RECT 1.722 1.096 1.733 1.225 ;
      RECT 2.528 1.068 2.574 1.196 ;
      RECT 1.676 1.068 1.722 1.196 ;
      RECT 3.232 0.655 3.322 1.23 ;
      RECT 2.49 1.121 2.623 1.154 ;
      RECT 2.11 1.121 2.243 1.154 ;
      RECT 2.194 1.05 2.205 1.179 ;
      RECT 1.638 1.121 1.771 1.154 ;
      RECT 1.161 1.121 1.294 1.154 ;
      RECT 1.245 1.05 1.256 1.179 ;
      RECT 0.69 0.465 0.78 1.23 ;
      RECT 2.205 1.045 2.528 1.135 ;
      RECT 1.256 1.045 1.676 1.135 ;
      RECT 2.148 1.079 2.194 1.207 ;
      RECT 1.199 1.079 1.245 1.207 ;
      RECT 0.045 0.96 0.78 1.05 ;
      RECT 0.045 0.252 0.135 1.05 ;
      RECT 0.045 0.252 0.185 0.342 ;
      RECT 2.652 0.71 2.742 0.991 ;
      RECT 2.652 0.71 2.858 0.8 ;
      RECT 2.768 0.35 2.858 0.8 ;
      RECT 1.255 0.505 2.037 0.595 ;
      RECT 1.947 0.35 2.037 0.595 ;
      RECT 1.947 0.35 2.858 0.44 ;
      RECT 1.87 0.685 2.01 0.855 ;
      RECT 1.05 0.685 2.45 0.775 ;
      RECT 2.36 0.53 2.45 0.775 ;
      RECT 1.05 0.325 1.14 0.775 ;
      RECT 2.36 0.53 2.678 0.62 ;
      RECT 1.05 0.325 1.857 0.415 ;
      RECT 1.767 0.205 1.857 0.415 ;
      RECT 1.809 0.96 2.071 1.05 ;
      RECT 1.798 0.916 1.809 1.045 ;
      RECT 0.87 0.245 0.96 1.03 ;
      RECT 1.798 0.96 2.117 1.027 ;
      RECT 1.752 0.888 1.798 1.016 ;
      RECT 2.033 0.941 2.166 0.974 ;
      RECT 2.117 0.87 2.128 0.999 ;
      RECT 1.714 0.941 1.847 0.974 ;
      RECT 2.128 0.865 2.33 0.955 ;
      RECT 0.87 0.865 1.752 0.955 ;
      RECT 2.071 0.899 2.33 0.955 ;
      RECT 0.805 0.245 0.96 0.335 ;
  END
END DFFSX1H7R

MACRO DFFSX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSX2H7R 0 0 ;
  SIZE 5.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.6 1.48 ;
        RECT 5.317 0.855 5.407 1.48 ;
        RECT 4.387 1.225 4.527 1.48 ;
        RECT 3.555 1.225 3.695 1.48 ;
        RECT 2.312 1.225 2.452 1.48 ;
        RECT 1.46 1.225 1.6 1.48 ;
        RECT 0.31 1.14 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.6 0.08 ;
        RECT 5.317 -0.08 5.407 0.353 ;
        RECT 4.807 -0.08 4.897 0.332 ;
        RECT 4.307 -0.08 4.397 0.33 ;
        RECT 3.802 -0.08 3.942 0.34 ;
        RECT 1.42 -0.08 1.56 0.175 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.425 0.345 0.65 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.6 0.545 0.87 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.067 0.21 5.157 1.146 ;
        RECT 5.035 0.21 5.157 0.375 ;
      LAYER MET2 ;
        RECT 5.05 0.18 5.15 0.56 ;
      LAYER VIA1 ;
        RECT 5.055 0.255 5.145 0.345 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.625 0.805 4.775 0.945 ;
        RECT 4.625 0.232 4.715 0.945 ;
        RECT 4.527 0.232 4.715 0.322 ;
      LAYER MET2 ;
        RECT 4.65 0.625 4.75 1.16 ;
      LAYER VIA1 ;
        RECT 4.655 0.855 4.745 0.945 ;
    END
  END QN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.65 0.625 3.785 0.825 ;
      LAYER MET2 ;
        RECT 3.65 0.43 3.75 0.96 ;
      LAYER VIA1 ;
        RECT 3.655 0.655 3.745 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 3.462 1.045 4.977 1.135 ;
      RECT 4.887 0.551 4.977 1.135 ;
      RECT 4.445 0.42 4.535 1.135 ;
      RECT 3.462 0.655 3.552 1.135 ;
      RECT 4.105 0.42 4.535 0.51 ;
      RECT 4.103 0.42 4.535 0.509 ;
      RECT 4.057 0.295 4.147 0.485 ;
      RECT 2.877 0.89 3.038 0.98 ;
      RECT 2.948 0.355 3.038 0.98 ;
      RECT 3.907 0.557 3.997 0.955 ;
      RECT 3.907 0.6 4.355 0.69 ;
      RECT 3.894 0.482 3.907 0.611 ;
      RECT 3.894 0.589 4.018 0.611 ;
      RECT 3.848 0.453 3.894 0.581 ;
      RECT 3.848 0.512 3.953 0.581 ;
      RECT 3.81 0.512 3.953 0.539 ;
      RECT 2.948 0.43 3.848 0.52 ;
      RECT 2.948 0.355 3.088 0.52 ;
      RECT 3.552 0.17 3.692 0.34 ;
      RECT 2.1 0.17 3.692 0.26 ;
      RECT 2.585 1.14 3.347 1.23 ;
      RECT 1.733 1.14 2.148 1.23 ;
      RECT 0.69 1.14 1.199 1.23 ;
      RECT 2.574 1.096 2.585 1.225 ;
      RECT 1.722 1.096 1.733 1.225 ;
      RECT 2.528 1.068 2.574 1.196 ;
      RECT 1.676 1.068 1.722 1.196 ;
      RECT 3.232 0.655 3.322 1.23 ;
      RECT 2.49 1.121 2.623 1.154 ;
      RECT 2.11 1.121 2.243 1.154 ;
      RECT 2.194 1.05 2.205 1.179 ;
      RECT 1.638 1.121 1.771 1.154 ;
      RECT 1.161 1.121 1.294 1.154 ;
      RECT 1.245 1.05 1.256 1.179 ;
      RECT 0.69 0.465 0.78 1.23 ;
      RECT 2.205 1.045 2.528 1.135 ;
      RECT 1.256 1.045 1.676 1.135 ;
      RECT 2.148 1.079 2.194 1.207 ;
      RECT 1.199 1.079 1.245 1.207 ;
      RECT 0.045 0.96 0.78 1.05 ;
      RECT 0.045 0.252 0.135 1.05 ;
      RECT 0.045 0.252 0.185 0.342 ;
      RECT 2.652 0.71 2.742 0.991 ;
      RECT 2.652 0.71 2.858 0.8 ;
      RECT 2.768 0.35 2.858 0.8 ;
      RECT 1.255 0.505 2.037 0.595 ;
      RECT 1.947 0.35 2.037 0.595 ;
      RECT 1.947 0.35 2.858 0.44 ;
      RECT 1.87 0.685 2.01 0.855 ;
      RECT 1.05 0.685 2.45 0.775 ;
      RECT 2.36 0.53 2.45 0.775 ;
      RECT 1.05 0.325 1.14 0.775 ;
      RECT 2.36 0.53 2.678 0.62 ;
      RECT 1.05 0.325 1.857 0.415 ;
      RECT 1.767 0.205 1.857 0.415 ;
      RECT 1.809 0.96 2.071 1.05 ;
      RECT 1.798 0.916 1.809 1.045 ;
      RECT 0.87 0.245 0.96 1.03 ;
      RECT 1.798 0.96 2.117 1.027 ;
      RECT 1.752 0.888 1.798 1.016 ;
      RECT 2.033 0.941 2.166 0.974 ;
      RECT 2.117 0.87 2.128 0.999 ;
      RECT 1.714 0.941 1.847 0.974 ;
      RECT 2.128 0.865 2.33 0.955 ;
      RECT 0.87 0.865 1.752 0.955 ;
      RECT 2.071 0.899 2.33 0.955 ;
      RECT 0.805 0.245 0.96 0.335 ;
  END
END DFFSX2H7R

MACRO DFFTRQX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFTRQX0P5H7R 0 0 ;
  SIZE 5.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.4 1.48 ;
        RECT 4.676 1.035 4.766 1.48 ;
        RECT 3.745 1.06 3.885 1.48 ;
        RECT 2.515 1.24 2.655 1.48 ;
        RECT 1.475 1.095 1.615 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.4 0.08 ;
        RECT 4.866 -0.08 4.956 0.33 ;
        RECT 3.836 -0.08 3.926 0.33 ;
        RECT 2.41 -0.08 2.55 0.305 ;
        RECT 1.505 -0.08 1.645 0.16 ;
        RECT 0.045 -0.08 0.185 0.32 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 4.606 0.643 4.781 0.869 ;
      LAYER MET2 ;
        RECT 4.65 0.425 4.75 0.96 ;
      LAYER VIA1 ;
        RECT 4.655 0.655 4.745 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.045 0.652 0.26 0.825 ;
        RECT 0.045 0.615 0.165 0.825 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.116 0.827 5.351 0.917 ;
        RECT 5.251 0.42 5.351 0.917 ;
        RECT 5.116 0.42 5.351 0.55 ;
        RECT 5.116 0.827 5.206 1.147 ;
        RECT 5.116 0.19 5.206 0.55 ;
      LAYER MET2 ;
        RECT 5.25 0.225 5.35 0.76 ;
      LAYER VIA1 ;
        RECT 5.255 0.455 5.345 0.545 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.375 0.41 0.49 0.645 ;
        RECT 0.224 0.41 0.49 0.545 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END RN
  OBS
    LAYER MET1 ;
      RECT 3.229 0.875 3.38 0.965 ;
      RECT 3.29 0.234 3.38 0.965 ;
      RECT 5.013 0.647 5.161 0.737 ;
      RECT 5.005 0.605 5.013 0.733 ;
      RECT 4.959 0.578 5.005 0.706 ;
      RECT 4.913 0.532 4.959 0.66 ;
      RECT 4.913 0.628 5.051 0.66 ;
      RECT 4.867 0.486 4.913 0.614 ;
      RECT 3.656 0.505 4.106 0.595 ;
      RECT 4.016 0.17 4.106 0.595 ;
      RECT 4.829 0.532 4.959 0.572 ;
      RECT 4.686 0.463 4.867 0.553 ;
      RECT 3.656 0.29 3.746 0.595 ;
      RECT 4.686 0.249 4.776 0.553 ;
      RECT 3.641 0.29 3.746 0.332 ;
      RECT 3.215 0.234 3.679 0.324 ;
      RECT 4.675 0.175 4.686 0.304 ;
      RECT 3.215 0.257 3.725 0.324 ;
      RECT 4.637 0.249 4.776 0.279 ;
      RECT 4.016 0.17 4.675 0.26 ;
      RECT 4.016 0.204 4.732 0.26 ;
      RECT 4.006 1.14 4.516 1.23 ;
      RECT 4.426 0.35 4.516 1.23 ;
      RECT 2.81 1.14 3.56 1.23 ;
      RECT 3.47 0.425 3.56 1.23 ;
      RECT 0.76 1.14 1.235 1.23 ;
      RECT 1.145 0.87 1.235 1.23 ;
      RECT 2.768 1.081 2.81 1.209 ;
      RECT 1.705 1.095 2.44 1.185 ;
      RECT 2.73 1.14 3.56 1.169 ;
      RECT 1.705 1.095 2.475 1.168 ;
      RECT 2.437 1.06 2.768 1.15 ;
      RECT 4.006 0.88 4.096 1.23 ;
      RECT 1.705 1.121 2.848 1.15 ;
      RECT 0.76 0.505 0.85 1.23 ;
      RECT 2.402 1.077 2.44 1.185 ;
      RECT 1.705 0.905 1.795 1.185 ;
      RECT 1.145 0.905 1.795 0.995 ;
      RECT 3.47 0.88 4.096 0.97 ;
      RECT 1.145 0.87 1.285 0.995 ;
      RECT 4.426 0.35 4.596 0.44 ;
      RECT 4.196 0.35 4.286 1.05 ;
      RECT 3.66 0.685 4.286 0.775 ;
      RECT 4.196 0.35 4.336 0.465 ;
      RECT 2.22 0.755 2.36 1.005 ;
      RECT 2.22 0.755 2.87 0.845 ;
      RECT 2.78 0.395 2.87 0.845 ;
      RECT 2.78 0.585 3.2 0.675 ;
      RECT 3.064 0.535 3.2 0.675 ;
      RECT 1.12 0.25 1.21 0.555 ;
      RECT 2.185 0.395 2.87 0.485 ;
      RECT 2.185 0.17 2.275 0.485 ;
      RECT 1.12 0.25 1.737 0.34 ;
      RECT 1.12 0.25 1.817 0.279 ;
      RECT 1.779 0.17 2.275 0.26 ;
      RECT 1.699 0.231 2.275 0.26 ;
      RECT 1.737 0.191 1.779 0.319 ;
      RECT 1.885 0.35 1.975 1.005 ;
      RECT 1.885 0.575 2.69 0.665 ;
      RECT 1.325 0.44 1.975 0.53 ;
      RECT 1.885 0.35 2.055 0.465 ;
      RECT 0.94 0.23 1.03 1.05 ;
      RECT 0.94 0.645 1.795 0.735 ;
      RECT 0.76 0.23 1.03 0.32 ;
      RECT 0.07 0.959 0.16 1.175 ;
      RECT 0.545 0.915 0.67 1.078 ;
      RECT 0.58 0.205 0.67 1.078 ;
      RECT 0.07 0.959 0.175 1.013 ;
      RECT 0.137 0.915 0.67 1.005 ;
      RECT 0.116 0.925 0.67 1.005 ;
      RECT 0.505 0.205 0.67 0.32 ;
  END
END DFFTRQX0P5H7R

MACRO DFFTRQX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFTRQX1H7R 0 0 ;
  SIZE 5.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.4 1.48 ;
        RECT 4.676 1.035 4.766 1.48 ;
        RECT 3.745 1.06 3.885 1.48 ;
        RECT 2.515 1.24 2.655 1.48 ;
        RECT 1.475 1.095 1.615 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.4 0.08 ;
        RECT 4.866 -0.08 4.956 0.33 ;
        RECT 3.836 -0.08 3.926 0.33 ;
        RECT 2.41 -0.08 2.55 0.305 ;
        RECT 1.505 -0.08 1.645 0.16 ;
        RECT 0.045 -0.08 0.185 0.32 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 4.606 0.643 4.776 0.869 ;
      LAYER MET2 ;
        RECT 4.65 0.425 4.75 0.96 ;
      LAYER VIA1 ;
        RECT 4.655 0.655 4.745 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.045 0.65 0.26 0.825 ;
        RECT 0.045 0.622 0.17 0.825 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.116 0.827 5.351 0.917 ;
        RECT 5.251 0.425 5.351 0.917 ;
        RECT 5.116 0.425 5.351 0.557 ;
        RECT 5.116 0.827 5.206 1.147 ;
        RECT 5.116 0.19 5.206 0.557 ;
      LAYER MET2 ;
        RECT 5.25 0.225 5.35 0.76 ;
      LAYER VIA1 ;
        RECT 5.255 0.455 5.345 0.545 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.375 0.41 0.49 0.645 ;
        RECT 0.219 0.41 0.49 0.545 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END RN
  OBS
    LAYER MET1 ;
      RECT 3.229 0.875 3.38 0.965 ;
      RECT 3.29 0.234 3.38 0.965 ;
      RECT 5.013 0.647 5.161 0.737 ;
      RECT 5.005 0.605 5.013 0.733 ;
      RECT 4.959 0.578 5.005 0.706 ;
      RECT 4.913 0.532 4.959 0.66 ;
      RECT 4.913 0.628 5.051 0.66 ;
      RECT 4.867 0.486 4.913 0.614 ;
      RECT 3.656 0.505 4.106 0.595 ;
      RECT 4.016 0.17 4.106 0.595 ;
      RECT 4.829 0.532 4.959 0.572 ;
      RECT 4.686 0.463 4.867 0.553 ;
      RECT 3.656 0.29 3.746 0.595 ;
      RECT 4.686 0.249 4.776 0.553 ;
      RECT 3.641 0.29 3.746 0.332 ;
      RECT 3.215 0.234 3.679 0.324 ;
      RECT 4.675 0.175 4.686 0.304 ;
      RECT 3.215 0.257 3.725 0.324 ;
      RECT 4.637 0.249 4.776 0.279 ;
      RECT 4.016 0.17 4.675 0.26 ;
      RECT 4.016 0.204 4.732 0.26 ;
      RECT 4.006 1.14 4.516 1.23 ;
      RECT 4.426 0.35 4.516 1.23 ;
      RECT 2.81 1.14 3.56 1.23 ;
      RECT 3.47 0.425 3.56 1.23 ;
      RECT 0.76 1.14 1.235 1.23 ;
      RECT 1.145 0.87 1.235 1.23 ;
      RECT 2.768 1.081 2.81 1.209 ;
      RECT 1.705 1.095 2.44 1.185 ;
      RECT 2.73 1.14 3.56 1.169 ;
      RECT 1.705 1.095 2.475 1.168 ;
      RECT 2.437 1.06 2.768 1.15 ;
      RECT 4.006 0.88 4.096 1.23 ;
      RECT 1.705 1.121 2.848 1.15 ;
      RECT 0.76 0.505 0.85 1.23 ;
      RECT 2.402 1.077 2.44 1.185 ;
      RECT 1.705 0.905 1.795 1.185 ;
      RECT 1.145 0.905 1.795 0.995 ;
      RECT 3.47 0.88 4.096 0.97 ;
      RECT 1.145 0.87 1.285 0.995 ;
      RECT 4.426 0.35 4.596 0.44 ;
      RECT 4.196 0.35 4.286 1.05 ;
      RECT 3.66 0.685 4.286 0.775 ;
      RECT 4.196 0.35 4.336 0.465 ;
      RECT 2.22 0.755 2.36 1.005 ;
      RECT 2.22 0.755 2.87 0.845 ;
      RECT 2.78 0.395 2.87 0.845 ;
      RECT 2.78 0.585 3.2 0.675 ;
      RECT 3.064 0.535 3.2 0.675 ;
      RECT 1.12 0.25 1.21 0.555 ;
      RECT 2.185 0.395 2.87 0.485 ;
      RECT 2.185 0.17 2.275 0.485 ;
      RECT 1.12 0.25 1.737 0.34 ;
      RECT 1.12 0.25 1.817 0.279 ;
      RECT 1.779 0.17 2.275 0.26 ;
      RECT 1.699 0.231 2.275 0.26 ;
      RECT 1.737 0.191 1.779 0.319 ;
      RECT 1.885 0.35 1.975 1.005 ;
      RECT 1.885 0.575 2.69 0.665 ;
      RECT 1.325 0.44 1.975 0.53 ;
      RECT 1.885 0.35 2.055 0.465 ;
      RECT 0.94 0.23 1.03 1.05 ;
      RECT 0.94 0.645 1.795 0.735 ;
      RECT 0.76 0.23 1.03 0.32 ;
      RECT 0.07 0.959 0.16 1.175 ;
      RECT 0.545 0.915 0.67 1.078 ;
      RECT 0.58 0.205 0.67 1.078 ;
      RECT 0.07 0.959 0.175 1.013 ;
      RECT 0.137 0.915 0.67 1.005 ;
      RECT 0.116 0.925 0.67 1.005 ;
      RECT 0.505 0.205 0.67 0.32 ;
  END
END DFFTRQX1H7R

MACRO DFFTRQX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFTRQX2H7R 0 0 ;
  SIZE 5.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.6 1.48 ;
        RECT 5.366 1.007 5.456 1.48 ;
        RECT 4.676 1.035 4.766 1.48 ;
        RECT 3.745 1.06 3.885 1.48 ;
        RECT 2.515 1.24 2.655 1.48 ;
        RECT 1.475 1.095 1.615 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.6 0.08 ;
        RECT 5.366 -0.08 5.456 0.33 ;
        RECT 4.866 -0.08 4.956 0.33 ;
        RECT 3.836 -0.08 3.926 0.33 ;
        RECT 2.41 -0.08 2.55 0.305 ;
        RECT 1.505 -0.08 1.645 0.16 ;
        RECT 0.045 -0.08 0.185 0.32 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 4.606 0.648 4.776 0.869 ;
      LAYER MET2 ;
        RECT 4.65 0.425 4.75 0.96 ;
      LAYER VIA1 ;
        RECT 4.655 0.655 4.745 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.045 0.637 0.26 0.825 ;
        RECT 0.045 0.605 0.155 0.825 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.116 0.827 5.417 0.917 ;
        RECT 5.327 0.435 5.417 0.917 ;
        RECT 5.116 0.435 5.417 0.545 ;
        RECT 5.116 0.827 5.206 1.147 ;
        RECT 5.116 0.19 5.206 0.545 ;
      LAYER MET2 ;
        RECT 5.25 0.225 5.35 0.76 ;
      LAYER VIA1 ;
        RECT 5.255 0.455 5.345 0.545 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.375 0.41 0.49 0.645 ;
        RECT 0.224 0.41 0.49 0.545 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END RN
  OBS
    LAYER MET1 ;
      RECT 3.229 0.875 3.38 0.965 ;
      RECT 3.29 0.234 3.38 0.965 ;
      RECT 5.013 0.647 5.237 0.737 ;
      RECT 5.005 0.605 5.013 0.733 ;
      RECT 4.959 0.578 5.005 0.706 ;
      RECT 4.913 0.532 4.959 0.66 ;
      RECT 4.913 0.628 5.051 0.66 ;
      RECT 4.867 0.486 4.913 0.614 ;
      RECT 3.656 0.505 4.106 0.595 ;
      RECT 4.016 0.17 4.106 0.595 ;
      RECT 4.829 0.532 4.959 0.572 ;
      RECT 4.686 0.463 4.867 0.553 ;
      RECT 3.656 0.29 3.746 0.595 ;
      RECT 4.686 0.249 4.776 0.553 ;
      RECT 3.641 0.29 3.746 0.332 ;
      RECT 3.215 0.234 3.679 0.324 ;
      RECT 4.675 0.175 4.686 0.304 ;
      RECT 3.215 0.257 3.725 0.324 ;
      RECT 4.637 0.249 4.776 0.279 ;
      RECT 4.016 0.17 4.675 0.26 ;
      RECT 4.016 0.204 4.732 0.26 ;
      RECT 4.006 1.14 4.516 1.23 ;
      RECT 4.426 0.35 4.516 1.23 ;
      RECT 2.81 1.14 3.56 1.23 ;
      RECT 3.47 0.425 3.56 1.23 ;
      RECT 0.76 1.14 1.235 1.23 ;
      RECT 1.145 0.87 1.235 1.23 ;
      RECT 2.768 1.081 2.81 1.209 ;
      RECT 1.705 1.095 2.44 1.185 ;
      RECT 2.73 1.14 3.56 1.169 ;
      RECT 1.705 1.095 2.475 1.168 ;
      RECT 2.437 1.06 2.768 1.15 ;
      RECT 4.006 0.88 4.096 1.23 ;
      RECT 1.705 1.121 2.848 1.15 ;
      RECT 0.76 0.505 0.85 1.23 ;
      RECT 2.402 1.077 2.44 1.185 ;
      RECT 1.705 0.905 1.795 1.185 ;
      RECT 1.145 0.905 1.795 0.995 ;
      RECT 3.47 0.88 4.096 0.97 ;
      RECT 1.145 0.87 1.285 0.995 ;
      RECT 4.426 0.35 4.596 0.44 ;
      RECT 4.196 0.35 4.286 1.05 ;
      RECT 3.66 0.685 4.286 0.775 ;
      RECT 4.196 0.35 4.336 0.465 ;
      RECT 2.22 0.755 2.36 1.005 ;
      RECT 2.22 0.755 2.87 0.845 ;
      RECT 2.78 0.395 2.87 0.845 ;
      RECT 2.78 0.585 3.2 0.675 ;
      RECT 3.064 0.535 3.2 0.675 ;
      RECT 1.12 0.25 1.21 0.555 ;
      RECT 2.185 0.395 2.87 0.485 ;
      RECT 2.185 0.17 2.275 0.485 ;
      RECT 1.12 0.25 1.737 0.34 ;
      RECT 1.12 0.25 1.817 0.279 ;
      RECT 1.779 0.17 2.275 0.26 ;
      RECT 1.699 0.231 2.275 0.26 ;
      RECT 1.737 0.191 1.779 0.319 ;
      RECT 1.885 0.35 1.975 1.005 ;
      RECT 1.885 0.575 2.69 0.665 ;
      RECT 1.325 0.44 1.975 0.53 ;
      RECT 1.885 0.35 2.055 0.465 ;
      RECT 0.94 0.23 1.03 1.05 ;
      RECT 0.94 0.645 1.795 0.735 ;
      RECT 0.76 0.23 1.03 0.32 ;
      RECT 0.07 0.959 0.16 1.175 ;
      RECT 0.545 0.915 0.67 1.078 ;
      RECT 0.58 0.205 0.67 1.078 ;
      RECT 0.07 0.959 0.175 1.013 ;
      RECT 0.137 0.915 0.67 1.005 ;
      RECT 0.116 0.925 0.67 1.005 ;
      RECT 0.505 0.205 0.67 0.32 ;
  END
END DFFTRQX2H7R

MACRO DFFX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFX0P5H7R 0 0 ;
  SIZE 4.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.6 1.48 ;
        RECT 4.094 1.19 4.234 1.48 ;
        RECT 3.319 1.19 3.459 1.48 ;
        RECT 2.286 1.225 2.426 1.48 ;
        RECT 1.455 1.14 1.595 1.48 ;
        RECT 0.31 1.11 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.6 0.08 ;
        RECT 4.119 -0.08 4.209 0.385 ;
        RECT 3.319 -0.08 3.459 0.21 ;
        RECT 2.288 -0.08 2.428 0.175 ;
        RECT 1.383 -0.08 1.523 0.185 ;
        RECT 0.32 -0.08 0.41 0.35 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.455 0.375 0.545 ;
        RECT 0.225 0.455 0.315 0.695 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.655 0.575 0.835 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.384 0.425 4.545 0.575 ;
        RECT 4.384 0.31 4.474 0.92 ;
      LAYER MET2 ;
        RECT 4.45 0.225 4.55 0.76 ;
      LAYER VIA1 ;
        RECT 4.455 0.455 4.545 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.455 0.795 3.739 0.885 ;
        RECT 3.455 0.3 3.724 0.39 ;
        RECT 3.455 0.3 3.545 0.885 ;
      LAYER MET2 ;
        RECT 3.45 0.225 3.55 0.76 ;
      LAYER VIA1 ;
        RECT 3.455 0.455 3.545 0.545 ;
    END
  END QN
  OBS
    LAYER MET1 ;
      RECT 2.843 1.075 3.156 1.165 ;
      RECT 2.843 1.075 3.174 1.156 ;
      RECT 2.843 1.075 3.216 1.126 ;
      RECT 3.174 0.267 3.221 1.103 ;
      RECT 4.094 0.595 4.184 1.1 ;
      RECT 3.118 1.056 4.184 1.1 ;
      RECT 3.174 1.01 4.184 1.1 ;
      RECT 3.156 1.028 4.184 1.1 ;
      RECT 3.174 0.291 3.264 1.1 ;
      RECT 2.777 0.265 3.216 0.355 ;
      RECT 3.854 0.31 3.944 0.92 ;
      RECT 3.749 0.585 3.944 0.675 ;
      RECT 1.99 1.14 2.132 1.23 ;
      RECT 1.99 1.14 2.178 1.207 ;
      RECT 2.094 1.121 2.224 1.161 ;
      RECT 2.132 1.079 2.224 1.161 ;
      RECT 2.178 1.033 2.27 1.115 ;
      RECT 2.224 0.987 2.316 1.069 ;
      RECT 2.27 0.941 2.359 1.025 ;
      RECT 2.27 0.941 2.397 0.984 ;
      RECT 2.994 0.465 3.084 0.965 ;
      RECT 2.316 0.896 3.084 0.965 ;
      RECT 2.359 0.875 3.084 0.965 ;
      RECT 1.05 0.302 1.14 0.575 ;
      RECT 2.705 0.465 3.084 0.555 ;
      RECT 2.691 0.42 2.705 0.548 ;
      RECT 2.645 0.39 2.691 0.518 ;
      RECT 2.599 0.344 2.645 0.472 ;
      RECT 2.599 0.446 2.743 0.472 ;
      RECT 2.553 0.298 2.599 0.426 ;
      RECT 1.05 0.302 1.577 0.392 ;
      RECT 2.515 0.344 2.645 0.384 ;
      RECT 1.05 0.302 1.623 0.369 ;
      RECT 2.048 0.275 2.553 0.365 ;
      RECT 1.539 0.283 1.669 0.323 ;
      RECT 1.577 0.241 1.671 0.299 ;
      RECT 1.577 0.241 1.709 0.279 ;
      RECT 2.048 0.17 2.138 0.365 ;
      RECT 1.671 0.17 2.138 0.26 ;
      RECT 1.623 0.195 2.138 0.26 ;
      RECT 1.669 0.171 1.671 0.299 ;
      RECT 0.68 1.14 1.216 1.23 ;
      RECT 1.126 0.875 1.216 1.23 ;
      RECT 0.68 0.46 0.77 1.23 ;
      RECT 1.126 0.96 1.997 1.05 ;
      RECT 1.126 0.96 2.043 1.027 ;
      RECT 0.045 0.93 0.77 1.02 ;
      RECT 1.076 0.875 1.216 0.965 ;
      RECT 1.959 0.941 2.089 0.981 ;
      RECT 2.089 0.813 2.123 0.941 ;
      RECT 1.997 0.899 2.123 0.941 ;
      RECT 2.043 0.853 2.089 0.981 ;
      RECT 0.045 0.275 0.135 1.02 ;
      RECT 2.123 0.695 2.169 0.901 ;
      RECT 2.123 0.695 2.213 0.856 ;
      RECT 2.123 0.695 2.803 0.785 ;
      RECT 0.045 0.275 0.185 0.365 ;
      RECT 1.41 0.78 1.915 0.87 ;
      RECT 1.825 0.35 1.915 0.87 ;
      RECT 1.41 0.72 1.5 0.87 ;
      RECT 1.825 0.515 2.533 0.605 ;
      RECT 1.753 0.35 1.915 0.44 ;
      RECT 0.87 0.265 0.96 1.045 ;
      RECT 0.87 0.695 1.32 0.785 ;
      RECT 1.23 0.51 1.32 0.785 ;
      RECT 1.23 0.51 1.694 0.6 ;
      RECT 0.805 0.265 0.96 0.355 ;
  END
END DFFX0P5H7R

MACRO DFFX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFX1H7R 0 0 ;
  SIZE 4.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.6 1.48 ;
        RECT 4.114 1.215 4.254 1.48 ;
        RECT 3.339 1.215 3.479 1.48 ;
        RECT 2.306 1.225 2.446 1.48 ;
        RECT 1.45 1.14 1.59 1.48 ;
        RECT 0.31 1.135 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.6 0.08 ;
        RECT 4.139 -0.08 4.229 0.365 ;
        RECT 3.359 -0.08 3.449 0.33 ;
        RECT 2.308 -0.08 2.448 0.23 ;
        RECT 1.36 -0.08 1.5 0.22 ;
        RECT 0.32 -0.08 0.41 0.35 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.455 0.375 0.545 ;
        RECT 0.225 0.455 0.315 0.695 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.595 0.555 0.865 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.379 0.805 4.545 0.895 ;
        RECT 4.455 0.335 4.545 0.895 ;
        RECT 4.379 0.335 4.545 0.425 ;
      LAYER MET2 ;
        RECT 4.45 0.225 4.55 0.76 ;
      LAYER VIA1 ;
        RECT 4.455 0.455 4.545 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.609 0.83 3.759 0.92 ;
        RECT 3.609 0.225 3.745 0.375 ;
        RECT 3.609 0.225 3.699 0.92 ;
      LAYER MET2 ;
        RECT 3.65 0.18 3.75 0.56 ;
      LAYER VIA1 ;
        RECT 3.655 0.255 3.745 0.345 ;
    END
  END QN
  OBS
    LAYER MET1 ;
      RECT 2.863 1.095 3.181 1.185 ;
      RECT 2.863 1.095 3.209 1.171 ;
      RECT 3.209 0.324 3.241 1.141 ;
      RECT 4.114 0.595 4.204 1.125 ;
      RECT 3.143 1.076 4.204 1.125 ;
      RECT 3.209 1.035 4.204 1.125 ;
      RECT 3.181 1.043 4.204 1.125 ;
      RECT 3.209 0.392 3.299 1.125 ;
      RECT 3.204 0.305 3.209 0.434 ;
      RECT 3.158 0.28 3.204 0.408 ;
      RECT 3.158 0.363 3.287 0.408 ;
      RECT 3.12 0.257 3.158 0.366 ;
      RECT 2.838 0.257 3.158 0.347 ;
      RECT 3.874 0.31 3.964 0.92 ;
      RECT 3.794 0.56 3.964 0.7 ;
      RECT 2.01 1.14 2.152 1.23 ;
      RECT 2.01 1.14 2.198 1.207 ;
      RECT 2.114 1.121 2.244 1.161 ;
      RECT 2.152 1.079 2.244 1.161 ;
      RECT 2.198 1.033 2.29 1.115 ;
      RECT 2.198 1.033 2.336 1.069 ;
      RECT 2.244 0.987 2.339 1.045 ;
      RECT 2.244 0.987 2.377 1.024 ;
      RECT 2.244 0.987 2.789 1.005 ;
      RECT 2.29 0.941 2.809 0.995 ;
      RECT 2.751 0.905 2.789 1.005 ;
      RECT 3.014 0.485 3.104 0.985 ;
      RECT 2.336 0.916 3.104 0.985 ;
      RECT 2.771 0.895 3.104 0.985 ;
      RECT 2.339 0.915 3.104 0.985 ;
      RECT 2.725 0.485 3.104 0.575 ;
      RECT 1.04 0.315 1.13 0.575 ;
      RECT 2.69 0.429 2.725 0.558 ;
      RECT 2.644 0.389 2.69 0.517 ;
      RECT 2.644 0.466 2.763 0.517 ;
      RECT 2.598 0.343 2.644 0.471 ;
      RECT 2.56 0.32 2.598 0.429 ;
      RECT 2.043 0.32 2.598 0.41 ;
      RECT 1.04 0.315 1.574 0.405 ;
      RECT 1.04 0.315 1.62 0.382 ;
      RECT 2.043 0.17 2.133 0.41 ;
      RECT 1.536 0.296 1.666 0.336 ;
      RECT 1.574 0.254 1.681 0.306 ;
      RECT 1.574 0.254 1.719 0.279 ;
      RECT 1.681 0.17 2.133 0.26 ;
      RECT 1.62 0.208 2.133 0.26 ;
      RECT 1.666 0.177 1.681 0.306 ;
      RECT 0.68 1.12 1.191 1.21 ;
      RECT 1.1 0.85 1.191 1.21 ;
      RECT 0.68 0.46 0.77 1.21 ;
      RECT 1.1 0.96 2.006 1.05 ;
      RECT 0.045 0.955 0.77 1.045 ;
      RECT 1.1 0.96 2.052 1.027 ;
      RECT 1.968 0.941 2.098 0.981 ;
      RECT 0.045 0.28 0.135 1.045 ;
      RECT 2.006 0.899 2.098 0.981 ;
      RECT 2.006 0.899 2.144 0.935 ;
      RECT 2.052 0.853 2.168 0.9 ;
      RECT 2.098 0.807 2.214 0.865 ;
      RECT 2.098 0.807 2.231 0.834 ;
      RECT 2.098 0.807 2.7 0.825 ;
      RECT 2.144 0.772 2.72 0.815 ;
      RECT 2.662 0.725 2.7 0.825 ;
      RECT 2.682 0.715 2.823 0.805 ;
      RECT 2.168 0.735 2.823 0.805 ;
      RECT 0.045 0.28 0.185 0.37 ;
      RECT 1.4 0.78 1.905 0.87 ;
      RECT 1.815 0.35 1.905 0.87 ;
      RECT 1.4 0.72 1.49 0.87 ;
      RECT 2.437 0.505 2.527 0.645 ;
      RECT 1.815 0.505 2.527 0.595 ;
      RECT 1.765 0.35 1.905 0.44 ;
      RECT 0.86 0.265 0.95 1.03 ;
      RECT 0.86 0.665 1.31 0.755 ;
      RECT 1.22 0.52 1.31 0.755 ;
      RECT 1.22 0.52 1.723 0.61 ;
      RECT 0.805 0.265 0.95 0.355 ;
  END
END DFFX1H7R

MACRO DFFX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFX2H7R 0 0 ;
  SIZE 5.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.6 1.48 ;
        RECT 5.325 0.93 5.415 1.48 ;
        RECT 4.785 1.225 4.925 1.48 ;
        RECT 4.29 1.225 4.43 1.48 ;
        RECT 3.73 1.225 3.87 1.48 ;
        RECT 2.475 1.225 2.615 1.48 ;
        RECT 1.98 1.225 2.12 1.48 ;
        RECT 1.42 1.225 1.56 1.48 ;
        RECT 0.295 1.075 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.6 0.08 ;
        RECT 5.325 -0.08 5.415 0.348 ;
        RECT 4.795 -0.08 4.885 0.345 ;
        RECT 4.27 -0.08 4.36 0.36 ;
        RECT 3.77 -0.08 3.86 0.38 ;
        RECT 2.56 -0.08 2.7 0.185 ;
        RECT 2.065 -0.08 2.205 0.185 ;
        RECT 1.37 -0.08 1.46 0.21 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.455 0.42 0.545 ;
        RECT 0.225 0.455 0.315 0.65 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.405 0.65 0.585 0.8 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.055 0.225 5.165 1.005 ;
      LAYER MET2 ;
        RECT 5.05 0.23 5.15 0.76 ;
      LAYER VIA1 ;
        RECT 5.055 0.455 5.145 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.01 0.855 4.175 0.955 ;
        RECT 4.01 0.24 4.11 0.955 ;
      LAYER MET2 ;
        RECT 4.05 0.63 4.15 1.16 ;
      LAYER VIA1 ;
        RECT 4.055 0.855 4.145 0.945 ;
    END
  END QN
  OBS
    LAYER MET1 ;
      RECT 3.184 1.095 3.538 1.185 ;
      RECT 3.184 1.095 3.555 1.177 ;
      RECT 3.555 0.323 3.588 1.152 ;
      RECT 4.725 0.591 4.815 1.135 ;
      RECT 3.5 1.076 4.815 1.135 ;
      RECT 3.555 1.045 4.815 1.135 ;
      RECT 3.538 1.048 4.815 1.135 ;
      RECT 3.555 0.391 3.645 1.135 ;
      RECT 3.513 0.286 3.555 0.414 ;
      RECT 3.513 0.363 3.634 0.414 ;
      RECT 3.475 0.265 3.513 0.374 ;
      RECT 3.285 0.265 3.513 0.355 ;
      RECT 4.545 0.31 4.635 0.92 ;
      RECT 4.355 0.585 4.635 0.675 ;
      RECT 2.21 1.045 2.922 1.135 ;
      RECT 3.11 0.895 3.465 0.985 ;
      RECT 3.375 0.48 3.465 0.985 ;
      RECT 2.924 0.48 3.465 0.57 ;
      RECT 1.07 0.302 1.497 0.392 ;
      RECT 2.027 0.275 2.681 0.365 ;
      RECT 1.07 0.17 1.16 0.392 ;
      RECT 1.667 0.17 1.884 0.26 ;
      RECT 0.97 0.17 1.16 0.26 ;
      RECT 3.072 0.895 3.11 1.004 ;
      RECT 3.052 0.905 3.072 1.033 ;
      RECT 3.006 0.938 3.052 1.066 ;
      RECT 2.96 0.984 3.006 1.112 ;
      RECT 2.922 1.026 2.96 1.135 ;
      RECT 2.886 0.461 2.924 0.57 ;
      RECT 2.857 0.427 2.886 0.556 ;
      RECT 2.811 0.39 2.857 0.518 ;
      RECT 2.765 0.344 2.811 0.472 ;
      RECT 2.719 0.298 2.765 0.426 ;
      RECT 2.681 0.275 2.719 0.384 ;
      RECT 1.989 0.256 2.027 0.365 ;
      RECT 1.968 0.226 1.989 0.355 ;
      RECT 1.922 0.193 1.968 0.321 ;
      RECT 1.884 0.17 1.922 0.279 ;
      RECT 1.629 0.17 1.667 0.279 ;
      RECT 1.627 0.171 1.629 0.299 ;
      RECT 1.581 0.195 1.627 0.323 ;
      RECT 1.535 0.241 1.581 0.369 ;
      RECT 1.497 0.283 1.535 0.392 ;
      RECT 0.68 1.12 1.16 1.21 ;
      RECT 1.07 0.85 1.16 1.21 ;
      RECT 1.935 0.85 2.025 1.135 ;
      RECT 1.07 1.045 2.025 1.135 ;
      RECT 0.68 0.44 0.77 1.21 ;
      RECT 0.045 0.89 0.77 0.98 ;
      RECT 1.935 0.85 2.831 0.94 ;
      RECT 1.935 0.85 2.877 0.917 ;
      RECT 0.045 0.28 0.135 0.98 ;
      RECT 2.793 0.831 2.923 0.871 ;
      RECT 2.11 0.673 2.2 0.94 ;
      RECT 2.831 0.789 2.933 0.843 ;
      RECT 2.831 0.789 2.971 0.819 ;
      RECT 2.933 0.71 3.201 0.8 ;
      RECT 2.877 0.743 3.201 0.8 ;
      RECT 2.923 0.715 2.933 0.843 ;
      RECT 0.045 0.28 0.185 0.37 ;
      RECT 1.33 0.865 1.845 0.955 ;
      RECT 1.755 0.35 1.845 0.955 ;
      RECT 1.33 0.815 1.42 0.955 ;
      RECT 2.665 0.577 2.755 0.76 ;
      RECT 2.636 0.494 2.665 0.623 ;
      RECT 2.598 0.532 2.711 0.589 ;
      RECT 1.755 0.48 2.636 0.57 ;
      RECT 1.705 0.35 1.845 0.44 ;
      RECT 0.86 0.538 0.95 1.03 ;
      RECT 0.86 0.538 1.665 0.628 ;
      RECT 0.89 0.35 0.98 0.628 ;
  END
END DFFX2H7R

MACRO DFFX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFX3H7R 0 0 ;
  SIZE 5.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.8 1.48 ;
        RECT 5.545 0.93 5.635 1.48 ;
        RECT 5.005 1.225 5.145 1.48 ;
        RECT 4.51 1.225 4.65 1.48 ;
        RECT 3.95 1.225 4.09 1.48 ;
        RECT 2.595 1.225 2.735 1.48 ;
        RECT 2.045 1.225 2.185 1.48 ;
        RECT 1.485 1.225 1.625 1.48 ;
        RECT 0.32 1.05 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.8 0.08 ;
        RECT 5.545 -0.08 5.635 0.363 ;
        RECT 5.015 -0.08 5.105 0.345 ;
        RECT 4.52 -0.08 4.61 0.35 ;
        RECT 4.005 -0.08 4.095 0.35 ;
        RECT 2.595 -0.08 2.735 0.21 ;
        RECT 2.099 -0.08 2.239 0.185 ;
        RECT 1.375 -0.08 1.515 0.185 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.455 0.375 0.545 ;
        RECT 0.225 0.455 0.315 0.695 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.405 0.635 0.605 0.77 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.295 0.295 5.385 0.905 ;
        RECT 5.255 0.425 5.385 0.575 ;
      LAYER MET2 ;
        RECT 5.25 0.225 5.35 0.76 ;
      LAYER VIA1 ;
        RECT 5.255 0.455 5.345 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.23 0.865 4.37 0.955 ;
        RECT 4.255 0.28 4.345 0.955 ;
      LAYER MET2 ;
        RECT 4.25 0.225 4.35 0.76 ;
      LAYER VIA1 ;
        RECT 4.255 0.455 4.345 0.545 ;
    END
  END QN
  OBS
    LAYER MET1 ;
      RECT 3.402 1.095 3.744 1.185 ;
      RECT 3.73 0.288 3.744 1.185 ;
      RECT 3.73 0.318 3.79 1.162 ;
      RECT 3.73 0.343 3.794 1.137 ;
      RECT 4.945 0.595 5.035 1.135 ;
      RECT 3.706 1.083 5.035 1.135 ;
      RECT 3.73 1.045 5.035 1.135 ;
      RECT 3.73 0.358 3.82 1.135 ;
      RECT 3.694 0.263 3.73 0.391 ;
      RECT 3.656 0.245 3.694 0.354 ;
      RECT 3.32 0.245 3.694 0.335 ;
      RECT 4.75 0.31 4.855 0.92 ;
      RECT 4.575 0.585 4.855 0.675 ;
      RECT 2.33 1.045 3.179 1.135 ;
      RECT 2.33 1.045 3.225 1.112 ;
      RECT 3.141 1.026 3.271 1.066 ;
      RECT 3.179 0.984 3.271 1.066 ;
      RECT 3.179 0.984 3.309 1.024 ;
      RECT 3.55 0.47 3.64 1.005 ;
      RECT 3.225 0.938 3.64 1.005 ;
      RECT 3.271 0.915 3.64 1.005 ;
      RECT 3.105 0.47 3.64 0.56 ;
      RECT 3.065 0.412 3.105 0.54 ;
      RECT 3.019 0.369 3.065 0.497 ;
      RECT 3.019 0.451 3.143 0.497 ;
      RECT 2.973 0.323 3.019 0.451 ;
      RECT 2.935 0.369 3.065 0.409 ;
      RECT 2.048 0.3 2.973 0.39 ;
      RECT 2.002 0.239 2.048 0.367 ;
      RECT 1.105 0.275 1.591 0.365 ;
      RECT 1.956 0.193 2.002 0.321 ;
      RECT 1.956 0.281 2.086 0.321 ;
      RECT 1.918 0.239 2.048 0.279 ;
      RECT 1.553 0.256 1.696 0.279 ;
      RECT 1.637 0.18 1.658 0.309 ;
      RECT 1.105 0.17 1.195 0.365 ;
      RECT 1.658 0.17 1.956 0.26 ;
      RECT 1 0.17 1.195 0.26 ;
      RECT 1.591 0.214 1.637 0.342 ;
      RECT 0.715 1.095 1.245 1.185 ;
      RECT 1.155 0.825 1.245 1.185 ;
      RECT 2.032 0.775 2.122 1.135 ;
      RECT 1.155 1.045 2.122 1.135 ;
      RECT 0.715 0.48 0.805 1.185 ;
      RECT 0.045 0.87 0.805 0.96 ;
      RECT 0.045 0.28 0.135 0.96 ;
      RECT 2.032 0.775 3.105 0.865 ;
      RECT 2.032 0.775 3.15 0.839 ;
      RECT 3.112 0.73 3.363 0.82 ;
      RECT 3.067 0.756 3.363 0.82 ;
      RECT 3.105 0.733 3.112 0.862 ;
      RECT 2.425 0.66 2.515 0.865 ;
      RECT 0.045 0.28 0.185 0.37 ;
      RECT 1.395 0.865 1.905 0.955 ;
      RECT 1.79 0.35 1.88 0.955 ;
      RECT 1.395 0.815 1.485 0.955 ;
      RECT 2.735 0.48 2.825 0.685 ;
      RECT 1.79 0.48 2.825 0.57 ;
      RECT 1.735 0.35 1.88 0.44 ;
      RECT 0.895 0.538 0.985 1.005 ;
      RECT 1.605 0.53 1.695 0.67 ;
      RECT 0.925 0.53 1.695 0.62 ;
      RECT 0.925 0.35 1.015 0.62 ;
  END
END DFFX3H7R

MACRO DLY1X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY1X2H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.1 0.855 1.19 1.48 ;
        RECT 0.33 1.07 0.42 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.06 -0.08 1.2 0.175 ;
        RECT 0.33 -0.08 0.42 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.775 0.385 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.35 1.025 1.545 1.175 ;
        RECT 1.35 0.265 1.44 1.175 ;
      LAYER MET2 ;
        RECT 1.45 0.84 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.82 0.665 0.91 1.075 ;
      RECT 0.82 0.665 1.26 0.755 ;
      RECT 1.17 0.265 1.26 0.755 ;
      RECT 0.82 0.265 1.26 0.365 ;
      RECT 0.82 0.225 0.91 0.365 ;
      RECT 0.59 0.205 0.68 1.155 ;
      RECT 0.59 0.46 1.035 0.55 ;
      RECT 0.07 0.205 0.16 1.155 ;
      RECT 0.41 0.445 0.5 0.585 ;
      RECT 0.07 0.445 0.5 0.535 ;
  END
END DLY1X2H7R

MACRO DLY1X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY1X6H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.59 0.87 1.68 1.48 ;
        RECT 1.09 0.855 1.18 1.48 ;
        RECT 0.33 1.07 0.42 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.59 -0.08 1.68 0.35 ;
        RECT 1.05 -0.08 1.19 0.175 ;
        RECT 0.33 -0.08 0.42 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.775 0.385 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.84 0.245 1.93 1.165 ;
        RECT 1.34 0.655 1.93 0.745 ;
        RECT 1.34 0.245 1.43 1.165 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.81 0.665 0.9 1.075 ;
      RECT 0.81 0.665 1.25 0.755 ;
      RECT 1.16 0.265 1.25 0.755 ;
      RECT 0.81 0.265 1.25 0.365 ;
      RECT 0.81 0.225 0.9 0.365 ;
      RECT 0.58 0.205 0.67 1.155 ;
      RECT 0.58 0.46 1.025 0.55 ;
      RECT 0.07 0.205 0.16 1.155 ;
      RECT 0.4 0.445 0.49 0.585 ;
      RECT 0.07 0.445 0.49 0.535 ;
  END
END DLY1X6H7R

MACRO DLY2X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY2X2H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.21 0.855 1.3 1.48 ;
        RECT 0.33 1.07 0.42 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.17 -0.08 1.31 0.175 ;
        RECT 0.33 -0.08 0.42 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.775 0.385 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.43 1.025 1.55 1.175 ;
        RECT 1.46 0.245 1.55 1.175 ;
      LAYER MET2 ;
        RECT 1.45 0.84 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.87 0.665 0.96 1.14 ;
      RECT 0.87 0.665 1.37 0.755 ;
      RECT 1.28 0.265 1.37 0.755 ;
      RECT 0.87 0.265 1.37 0.365 ;
      RECT 0.87 0.225 0.96 0.365 ;
      RECT 0.64 0.205 0.73 1.155 ;
      RECT 0.64 0.46 1.145 0.55 ;
      RECT 0.07 0.205 0.16 1.155 ;
      RECT 0.07 0.47 0.55 0.56 ;
  END
END DLY2X2H7R

MACRO DLY2X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY2X6H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.71 0.87 1.8 1.48 ;
        RECT 1.21 0.855 1.3 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.71 -0.08 1.8 0.35 ;
        RECT 1.17 -0.08 1.31 0.175 ;
        RECT 0.33 -0.08 0.42 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.775 0.385 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.96 0.245 2.05 1.165 ;
        RECT 1.46 0.655 2.05 0.745 ;
        RECT 1.46 0.245 1.55 1.155 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.87 0.665 0.96 1.085 ;
      RECT 0.87 0.665 1.37 0.755 ;
      RECT 1.28 0.265 1.37 0.755 ;
      RECT 0.87 0.265 1.37 0.365 ;
      RECT 0.87 0.225 0.96 0.365 ;
      RECT 0.64 0.205 0.73 1.155 ;
      RECT 0.64 0.46 1.145 0.55 ;
      RECT 0.07 0.205 0.16 1.155 ;
      RECT 0.07 0.47 0.55 0.56 ;
  END
END DLY2X6H7R

MACRO DLY3X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY3X2H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.35 0.855 1.44 1.48 ;
        RECT 0.33 1.07 0.42 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.29 -0.08 1.43 0.175 ;
        RECT 0.33 -0.08 0.42 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.775 0.385 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.6 1.025 1.745 1.175 ;
        RECT 1.6 0.245 1.69 1.175 ;
      LAYER MET2 ;
        RECT 1.65 0.84 1.75 1.22 ;
      LAYER VIA1 ;
        RECT 1.655 1.055 1.745 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.93 0.665 1.02 1.145 ;
      RECT 0.93 0.665 1.47 0.755 ;
      RECT 1.38 0.265 1.47 0.755 ;
      RECT 0.93 0.265 1.47 0.365 ;
      RECT 0.93 0.225 1.02 0.365 ;
      RECT 0.7 0.205 0.79 1.155 ;
      RECT 0.7 0.46 1.145 0.55 ;
      RECT 0.07 0.205 0.16 1.155 ;
      RECT 0.07 0.47 0.55 0.56 ;
  END
END DLY3X2H7R

MACRO DLY3X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY3X6H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 1.85 1.07 1.94 1.48 ;
        RECT 1.35 0.855 1.44 1.48 ;
        RECT 0.33 1.07 0.42 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 1.825 -0.08 1.965 0.325 ;
        RECT 1.29 -0.08 1.43 0.175 ;
        RECT 0.33 -0.08 0.42 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.775 0.385 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.1 0.245 2.19 1.175 ;
        RECT 1.6 0.855 2.19 0.945 ;
        RECT 1.6 0.415 2.19 0.505 ;
        RECT 1.6 0.855 1.69 1.195 ;
        RECT 1.6 0.28 1.69 0.505 ;
      LAYER MET2 ;
        RECT 2.05 0.63 2.15 1.16 ;
      LAYER VIA1 ;
        RECT 2.055 0.855 2.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.93 0.665 1.02 1.145 ;
      RECT 0.93 0.665 1.355 0.755 ;
      RECT 1.265 0.265 1.355 0.755 ;
      RECT 1.265 0.6 1.925 0.69 ;
      RECT 0.93 0.265 1.355 0.365 ;
      RECT 0.93 0.225 1.02 0.365 ;
      RECT 0.7 0.205 0.79 1.155 ;
      RECT 0.7 0.47 1.175 0.56 ;
      RECT 0.07 0.205 0.16 1.155 ;
      RECT 0.07 0.47 0.595 0.56 ;
  END
END DLY3X6H7R

MACRO DLY4X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY4X2H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.435 1.069 1.525 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.41 -0.08 1.55 0.37 ;
        RECT 0.295 -0.08 0.435 0.37 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.575 0.39 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.655 1.025 1.807 1.175 ;
        RECT 1.717 0.295 1.807 1.175 ;
        RECT 1.66 0.295 1.807 0.385 ;
      LAYER MET2 ;
        RECT 1.65 0.84 1.75 1.22 ;
      LAYER VIA1 ;
        RECT 1.655 1.055 1.745 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.005 0.84 1.095 1.155 ;
      RECT 1.005 0.84 1.616 0.93 ;
      RECT 1.526 0.48 1.616 0.93 ;
      RECT 1.005 0.48 1.616 0.57 ;
      RECT 1.005 0.27 1.095 0.57 ;
      RECT 0.775 0.27 0.865 1.177 ;
      RECT 0.775 0.66 1.27 0.75 ;
      RECT 0.07 0.27 0.16 1.155 ;
      RECT 0.07 0.88 0.649 0.97 ;
      RECT 0.559 0.63 0.649 0.97 ;
  END
END DLY4X2H7R

MACRO DLY4X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY4X6H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 2.035 1.07 2.125 1.48 ;
        RECT 1.435 1.07 1.525 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 2.035 -0.08 2.125 0.396 ;
        RECT 1.41 -0.08 1.55 0.37 ;
        RECT 0.32 -0.08 0.41 0.37 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.575 0.39 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.285 0.31 2.375 0.965 ;
        RECT 1.855 0.874 2.375 0.965 ;
        RECT 1.748 0.956 1.945 1.046 ;
        RECT 1.855 0.32 1.945 1.046 ;
        RECT 1.748 0.32 1.945 0.41 ;
      LAYER MET2 ;
        RECT 1.85 0.225 1.95 0.76 ;
      LAYER VIA1 ;
        RECT 1.855 0.455 1.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.005 0.82 1.095 1.125 ;
      RECT 1.005 0.82 1.669 0.91 ;
      RECT 1.579 0.46 1.669 0.91 ;
      RECT 1.579 0.615 1.763 0.755 ;
      RECT 1.005 0.46 1.669 0.55 ;
      RECT 1.005 0.27 1.095 0.55 ;
      RECT 0.775 0.245 0.865 1.157 ;
      RECT 0.775 0.64 1.27 0.73 ;
      RECT 0.07 0.245 0.16 1.155 ;
      RECT 0.07 0.88 0.649 0.97 ;
      RECT 0.559 0.43 0.649 0.97 ;
  END
END DLY4X6H7R

MACRO EDFFQX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFQX0P5H7R 0 0 ;
  SIZE 7 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7 1.48 ;
        RECT 6.552 0.855 6.642 1.48 ;
        RECT 6.161 1.225 6.301 1.48 ;
        RECT 4.799 1.225 4.939 1.48 ;
        RECT 3.087 1.24 3.227 1.48 ;
        RECT 1.522 1.225 1.662 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7 0.08 ;
        RECT 6.249 -0.08 6.389 0.305 ;
        RECT 5.656 -0.08 5.796 0.305 ;
        RECT 4.989 -0.08 5.079 0.366 ;
        RECT 4.339 -0.08 4.429 0.39 ;
        RECT 3.174 -0.08 3.314 0.175 ;
        RECT 1.537 -0.08 1.681 0.355 ;
        RECT 0.295 -0.08 0.435 0.339 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.625 0.45 1.79 0.651 ;
      LAYER MET2 ;
        RECT 1.65 0.23 1.75 0.76 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.625 0.608 0.818 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.568 1.14 1.099 1.23 ;
        RECT 0.568 0.915 0.658 1.23 ;
        RECT 0.25 0.915 0.658 1.005 ;
        RECT 0.25 0.644 0.35 1.005 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.802 0.65 6.892 1.039 ;
        RECT 6.53 0.65 6.892 0.75 ;
        RECT 6.53 0.186 6.62 0.75 ;
      LAYER MET2 ;
        RECT 6.65 0.425 6.75 0.96 ;
      LAYER VIA1 ;
        RECT 6.655 0.655 6.745 0.745 ;
    END
  END Q
  OBS
    LAYER MET1 ;
      RECT 5.11 1.14 5.99 1.23 ;
      RECT 3.384 1.14 4.331 1.23 ;
      RECT 1.833 1.14 2.87 1.23 ;
      RECT 1.249 1.14 1.351 1.23 ;
      RECT 2.988 1.06 3.266 1.15 ;
      RECT 4.464 1.045 4.977 1.135 ;
      RECT 1.484 1.045 1.7 1.135 ;
      RECT 6.174 0.994 6.385 1.084 ;
      RECT 6.295 0.853 6.385 1.084 ;
      RECT 6.35 0.399 6.44 0.943 ;
      RECT 5.77 0.399 6.44 0.489 ;
      RECT 6.024 0.205 6.114 0.489 ;
      RECT 6.136 0.994 6.174 1.103 ;
      RECT 6.12 1.002 6.136 1.13 ;
      RECT 6.074 1.033 6.12 1.161 ;
      RECT 6.028 1.079 6.074 1.207 ;
      RECT 5.99 1.121 6.028 1.23 ;
      RECT 5.072 1.121 5.11 1.23 ;
      RECT 5.061 1.096 5.072 1.225 ;
      RECT 5.015 1.068 5.061 1.196 ;
      RECT 4.977 1.045 5.015 1.154 ;
      RECT 4.426 1.045 4.464 1.154 ;
      RECT 4.415 1.05 4.426 1.179 ;
      RECT 4.369 1.079 4.415 1.207 ;
      RECT 4.331 1.121 4.369 1.23 ;
      RECT 3.346 1.121 3.384 1.23 ;
      RECT 3.304 1.081 3.346 1.209 ;
      RECT 3.266 1.06 3.304 1.169 ;
      RECT 2.95 1.06 2.988 1.169 ;
      RECT 2.908 1.081 2.95 1.209 ;
      RECT 2.87 1.121 2.908 1.23 ;
      RECT 1.795 1.121 1.833 1.23 ;
      RECT 1.784 1.096 1.795 1.225 ;
      RECT 1.738 1.068 1.784 1.196 ;
      RECT 1.7 1.045 1.738 1.154 ;
      RECT 1.446 1.045 1.484 1.154 ;
      RECT 1.435 1.05 1.446 1.179 ;
      RECT 1.389 1.079 1.435 1.207 ;
      RECT 1.351 1.121 1.389 1.23 ;
      RECT 5.148 0.96 5.808 1.05 ;
      RECT 5.137 0.916 5.148 1.045 ;
      RECT 5.137 0.96 5.854 1.027 ;
      RECT 5.091 0.888 5.137 1.016 ;
      RECT 4.039 0.806 4.129 0.987 ;
      RECT 5.77 0.941 5.889 0.987 ;
      RECT 5.053 0.941 5.186 0.974 ;
      RECT 4.039 0.865 5.091 0.955 ;
      RECT 5.808 0.899 5.935 0.946 ;
      RECT 5.854 0.858 5.889 0.987 ;
      RECT 5.889 0.579 5.979 0.901 ;
      RECT 4.025 0.731 4.039 0.859 ;
      RECT 3.981 0.761 4.085 0.83 ;
      RECT 3.935 0.35 4.025 0.785 ;
      RECT 6.119 0.579 6.26 0.71 ;
      RECT 5.406 0.579 6.26 0.669 ;
      RECT 5.406 0.23 5.496 0.669 ;
      RECT 3.854 0.35 4.025 0.44 ;
      RECT 5.194 0.23 5.496 0.32 ;
      RECT 5.226 0.78 5.695 0.87 ;
      RECT 5.555 0.759 5.695 0.87 ;
      RECT 2.359 0.17 2.449 0.82 ;
      RECT 5.226 0.481 5.316 0.87 ;
      RECT 4.115 0.481 5.316 0.571 ;
      RECT 4.735 0.266 4.825 0.571 ;
      RECT 4.115 0.17 4.205 0.571 ;
      RECT 3.086 0.265 3.39 0.355 ;
      RECT 3.075 0.221 3.086 0.35 ;
      RECT 3.075 0.265 3.436 0.332 ;
      RECT 3.029 0.193 3.075 0.321 ;
      RECT 3.352 0.246 3.485 0.279 ;
      RECT 3.436 0.175 3.447 0.304 ;
      RECT 2.991 0.246 3.124 0.279 ;
      RECT 3.447 0.17 4.205 0.26 ;
      RECT 2.359 0.17 3.029 0.26 ;
      RECT 3.39 0.204 4.205 0.26 ;
      RECT 3.422 0.96 3.842 1.05 ;
      RECT 3.38 0.901 3.422 1.029 ;
      RECT 3.342 0.96 3.842 0.989 ;
      RECT 2.72 0.88 3.38 0.97 ;
      RECT 2.72 0.941 3.46 0.97 ;
      RECT 2.72 0.739 2.81 0.97 ;
      RECT 3.503 0.7 3.667 0.87 ;
      RECT 3.565 0.36 3.667 0.87 ;
      RECT 2.999 0.7 3.667 0.79 ;
      RECT 3.515 0.36 3.667 0.45 ;
      RECT 2.467 0.959 2.629 1.049 ;
      RECT 2.539 0.35 2.629 1.049 ;
      RECT 3.206 0.52 3.419 0.61 ;
      RECT 2.539 0.445 3.296 0.535 ;
      RECT 2.539 0.35 2.679 0.535 ;
      RECT 1.872 0.96 2.357 1.05 ;
      RECT 1.861 0.916 1.872 1.045 ;
      RECT 0.761 0.935 1.1 1.025 ;
      RECT 1.815 0.888 1.861 1.016 ;
      RECT 2.179 0.248 2.269 1.05 ;
      RECT 1.777 0.941 1.91 0.974 ;
      RECT 1.01 0.865 1.815 0.955 ;
      RECT 1.349 0.325 1.439 0.955 ;
      RECT 1.034 0.325 1.439 0.415 ;
      RECT 1.949 0.78 2.089 0.87 ;
      RECT 1.949 0.27 2.039 0.87 ;
      RECT 1.787 0.27 2.039 0.36 ;
      RECT 0.07 0.201 0.16 1.065 ;
      RECT 0.71 0.445 0.8 0.727 ;
      RECT 0.71 0.561 1.255 0.651 ;
      RECT 0.07 0.445 0.8 0.535 ;
      RECT 4.334 0.661 5.061 0.751 ;
  END
END EDFFQX0P5H7R

MACRO EDFFQX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFQX1H7R 0 0 ;
  SIZE 7 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7 1.48 ;
        RECT 6.552 0.855 6.642 1.48 ;
        RECT 6.161 1.225 6.301 1.48 ;
        RECT 4.799 1.225 4.939 1.48 ;
        RECT 3.087 1.24 3.227 1.48 ;
        RECT 1.522 1.225 1.662 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7 0.08 ;
        RECT 6.249 -0.08 6.389 0.305 ;
        RECT 5.656 -0.08 5.796 0.305 ;
        RECT 4.989 -0.08 5.079 0.366 ;
        RECT 4.339 -0.08 4.429 0.365 ;
        RECT 3.174 -0.08 3.314 0.175 ;
        RECT 1.537 -0.08 1.681 0.355 ;
        RECT 0.295 -0.08 0.435 0.339 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.625 0.45 1.777 0.651 ;
      LAYER MET2 ;
        RECT 1.65 0.23 1.75 0.76 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.625 0.608 0.818 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.568 1.14 1.099 1.23 ;
        RECT 0.568 0.915 0.658 1.23 ;
        RECT 0.25 0.915 0.658 1.005 ;
        RECT 0.25 0.644 0.35 1.005 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.802 0.65 6.892 1.099 ;
        RECT 6.53 0.65 6.892 0.75 ;
        RECT 6.53 0.186 6.62 0.75 ;
      LAYER MET2 ;
        RECT 6.65 0.425 6.75 0.96 ;
      LAYER VIA1 ;
        RECT 6.655 0.655 6.745 0.745 ;
    END
  END Q
  OBS
    LAYER MET1 ;
      RECT 5.11 1.14 5.99 1.23 ;
      RECT 3.384 1.14 4.331 1.23 ;
      RECT 1.833 1.14 2.87 1.23 ;
      RECT 1.249 1.14 1.351 1.23 ;
      RECT 2.988 1.06 3.266 1.15 ;
      RECT 4.464 1.045 4.977 1.135 ;
      RECT 1.484 1.045 1.7 1.135 ;
      RECT 6.174 0.994 6.385 1.084 ;
      RECT 6.295 0.853 6.385 1.084 ;
      RECT 6.35 0.399 6.44 0.943 ;
      RECT 5.77 0.399 6.44 0.489 ;
      RECT 6.024 0.205 6.114 0.489 ;
      RECT 6.136 0.994 6.174 1.103 ;
      RECT 6.12 1.002 6.136 1.13 ;
      RECT 6.074 1.033 6.12 1.161 ;
      RECT 6.028 1.079 6.074 1.207 ;
      RECT 5.99 1.121 6.028 1.23 ;
      RECT 5.072 1.121 5.11 1.23 ;
      RECT 5.061 1.096 5.072 1.225 ;
      RECT 5.015 1.068 5.061 1.196 ;
      RECT 4.977 1.045 5.015 1.154 ;
      RECT 4.426 1.045 4.464 1.154 ;
      RECT 4.415 1.05 4.426 1.179 ;
      RECT 4.369 1.079 4.415 1.207 ;
      RECT 4.331 1.121 4.369 1.23 ;
      RECT 3.346 1.121 3.384 1.23 ;
      RECT 3.304 1.081 3.346 1.209 ;
      RECT 3.266 1.06 3.304 1.169 ;
      RECT 2.95 1.06 2.988 1.169 ;
      RECT 2.908 1.081 2.95 1.209 ;
      RECT 2.87 1.121 2.908 1.23 ;
      RECT 1.795 1.121 1.833 1.23 ;
      RECT 1.784 1.096 1.795 1.225 ;
      RECT 1.738 1.068 1.784 1.196 ;
      RECT 1.7 1.045 1.738 1.154 ;
      RECT 1.446 1.045 1.484 1.154 ;
      RECT 1.435 1.05 1.446 1.179 ;
      RECT 1.389 1.079 1.435 1.207 ;
      RECT 1.351 1.121 1.389 1.23 ;
      RECT 5.148 0.96 5.808 1.05 ;
      RECT 5.137 0.916 5.148 1.045 ;
      RECT 5.137 0.96 5.854 1.027 ;
      RECT 5.091 0.888 5.137 1.016 ;
      RECT 4.039 0.806 4.129 0.987 ;
      RECT 5.77 0.941 5.889 0.987 ;
      RECT 5.053 0.941 5.186 0.974 ;
      RECT 4.039 0.865 5.091 0.955 ;
      RECT 5.808 0.899 5.935 0.946 ;
      RECT 5.854 0.858 5.889 0.987 ;
      RECT 5.889 0.579 5.979 0.901 ;
      RECT 4.025 0.731 4.039 0.859 ;
      RECT 3.981 0.761 4.085 0.83 ;
      RECT 3.935 0.35 4.025 0.785 ;
      RECT 6.119 0.579 6.26 0.71 ;
      RECT 5.406 0.579 6.26 0.669 ;
      RECT 5.406 0.23 5.496 0.669 ;
      RECT 3.854 0.35 4.025 0.44 ;
      RECT 5.194 0.23 5.496 0.32 ;
      RECT 5.226 0.78 5.695 0.87 ;
      RECT 5.555 0.759 5.695 0.87 ;
      RECT 2.359 0.17 2.449 0.82 ;
      RECT 5.226 0.456 5.316 0.87 ;
      RECT 4.115 0.456 5.316 0.546 ;
      RECT 4.735 0.266 4.825 0.546 ;
      RECT 4.115 0.17 4.205 0.546 ;
      RECT 3.086 0.265 3.39 0.355 ;
      RECT 3.075 0.221 3.086 0.35 ;
      RECT 3.075 0.265 3.436 0.332 ;
      RECT 3.029 0.193 3.075 0.321 ;
      RECT 3.352 0.246 3.485 0.279 ;
      RECT 3.436 0.175 3.447 0.304 ;
      RECT 2.991 0.246 3.124 0.279 ;
      RECT 3.447 0.17 4.205 0.26 ;
      RECT 2.359 0.17 3.029 0.26 ;
      RECT 3.39 0.204 4.205 0.26 ;
      RECT 3.422 0.96 3.842 1.05 ;
      RECT 3.38 0.901 3.422 1.029 ;
      RECT 3.342 0.96 3.842 0.989 ;
      RECT 2.72 0.88 3.38 0.97 ;
      RECT 2.72 0.941 3.46 0.97 ;
      RECT 2.72 0.739 2.81 0.97 ;
      RECT 3.503 0.7 3.667 0.87 ;
      RECT 3.565 0.36 3.667 0.87 ;
      RECT 2.999 0.7 3.667 0.79 ;
      RECT 3.515 0.36 3.667 0.45 ;
      RECT 2.467 0.959 2.629 1.049 ;
      RECT 2.539 0.35 2.629 1.049 ;
      RECT 3.206 0.52 3.419 0.61 ;
      RECT 2.539 0.445 3.296 0.535 ;
      RECT 2.539 0.35 2.679 0.535 ;
      RECT 1.872 0.96 2.357 1.05 ;
      RECT 1.861 0.916 1.872 1.045 ;
      RECT 0.761 0.935 1.1 1.025 ;
      RECT 1.815 0.888 1.861 1.016 ;
      RECT 2.179 0.228 2.269 1.05 ;
      RECT 1.777 0.941 1.91 0.974 ;
      RECT 1.01 0.865 1.815 0.955 ;
      RECT 1.349 0.325 1.439 0.955 ;
      RECT 1.034 0.325 1.439 0.415 ;
      RECT 1.949 0.78 2.089 0.87 ;
      RECT 1.949 0.27 2.039 0.87 ;
      RECT 1.787 0.27 2.039 0.36 ;
      RECT 0.07 0.201 0.16 1.065 ;
      RECT 0.71 0.445 0.8 0.727 ;
      RECT 0.71 0.561 1.255 0.651 ;
      RECT 0.07 0.445 0.8 0.535 ;
      RECT 4.334 0.661 5.061 0.751 ;
  END
END EDFFQX1H7R

MACRO EDFFQX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFQX2H7R 0 0 ;
  SIZE 7 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7 1.48 ;
        RECT 6.552 0.855 6.642 1.48 ;
        RECT 6.161 1.225 6.301 1.48 ;
        RECT 4.799 1.225 4.939 1.48 ;
        RECT 3.087 1.24 3.227 1.48 ;
        RECT 1.522 1.225 1.662 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7 0.08 ;
        RECT 6.78 -0.08 6.87 0.335 ;
        RECT 6.249 -0.08 6.389 0.305 ;
        RECT 5.656 -0.08 5.796 0.305 ;
        RECT 4.989 -0.08 5.079 0.366 ;
        RECT 4.339 -0.08 4.429 0.364 ;
        RECT 3.174 -0.08 3.314 0.175 ;
        RECT 1.537 -0.08 1.681 0.355 ;
        RECT 0.295 -0.08 0.435 0.339 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.625 0.45 1.777 0.651 ;
      LAYER MET2 ;
        RECT 1.65 0.23 1.75 0.76 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.625 0.608 0.818 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.568 1.14 1.099 1.23 ;
        RECT 0.568 0.915 0.658 1.23 ;
        RECT 0.25 0.915 0.658 1.005 ;
        RECT 0.25 0.644 0.35 1.005 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.802 0.65 6.892 1.099 ;
        RECT 6.53 0.65 6.892 0.75 ;
        RECT 6.53 0.186 6.62 0.75 ;
      LAYER MET2 ;
        RECT 6.65 0.425 6.75 0.96 ;
      LAYER VIA1 ;
        RECT 6.655 0.655 6.745 0.745 ;
    END
  END Q
  OBS
    LAYER MET1 ;
      RECT 5.11 1.14 5.99 1.23 ;
      RECT 3.384 1.14 4.331 1.23 ;
      RECT 1.833 1.14 2.87 1.23 ;
      RECT 1.249 1.14 1.351 1.23 ;
      RECT 2.988 1.06 3.266 1.15 ;
      RECT 4.464 1.045 4.977 1.135 ;
      RECT 1.484 1.045 1.7 1.135 ;
      RECT 6.174 0.994 6.385 1.084 ;
      RECT 6.295 0.853 6.385 1.084 ;
      RECT 6.35 0.399 6.44 0.943 ;
      RECT 5.77 0.399 6.44 0.489 ;
      RECT 6.024 0.205 6.114 0.489 ;
      RECT 6.136 0.994 6.174 1.103 ;
      RECT 6.12 1.002 6.136 1.13 ;
      RECT 6.074 1.033 6.12 1.161 ;
      RECT 6.028 1.079 6.074 1.207 ;
      RECT 5.99 1.121 6.028 1.23 ;
      RECT 5.072 1.121 5.11 1.23 ;
      RECT 5.061 1.096 5.072 1.225 ;
      RECT 5.015 1.068 5.061 1.196 ;
      RECT 4.977 1.045 5.015 1.154 ;
      RECT 4.426 1.045 4.464 1.154 ;
      RECT 4.415 1.05 4.426 1.179 ;
      RECT 4.369 1.079 4.415 1.207 ;
      RECT 4.331 1.121 4.369 1.23 ;
      RECT 3.346 1.121 3.384 1.23 ;
      RECT 3.304 1.081 3.346 1.209 ;
      RECT 3.266 1.06 3.304 1.169 ;
      RECT 2.95 1.06 2.988 1.169 ;
      RECT 2.908 1.081 2.95 1.209 ;
      RECT 2.87 1.121 2.908 1.23 ;
      RECT 1.795 1.121 1.833 1.23 ;
      RECT 1.784 1.096 1.795 1.225 ;
      RECT 1.738 1.068 1.784 1.196 ;
      RECT 1.7 1.045 1.738 1.154 ;
      RECT 1.446 1.045 1.484 1.154 ;
      RECT 1.435 1.05 1.446 1.179 ;
      RECT 1.389 1.079 1.435 1.207 ;
      RECT 1.351 1.121 1.389 1.23 ;
      RECT 5.148 0.96 5.808 1.05 ;
      RECT 5.137 0.916 5.148 1.045 ;
      RECT 5.137 0.96 5.854 1.027 ;
      RECT 5.091 0.888 5.137 1.016 ;
      RECT 4.039 0.806 4.129 0.987 ;
      RECT 5.77 0.941 5.889 0.987 ;
      RECT 5.053 0.941 5.186 0.974 ;
      RECT 4.039 0.865 5.091 0.955 ;
      RECT 5.808 0.899 5.935 0.946 ;
      RECT 5.854 0.858 5.889 0.987 ;
      RECT 5.889 0.579 5.979 0.901 ;
      RECT 4.025 0.731 4.039 0.859 ;
      RECT 3.981 0.761 4.085 0.83 ;
      RECT 3.935 0.35 4.025 0.785 ;
      RECT 6.119 0.579 6.26 0.71 ;
      RECT 5.406 0.579 6.26 0.669 ;
      RECT 5.406 0.23 5.496 0.669 ;
      RECT 3.854 0.35 4.025 0.44 ;
      RECT 5.194 0.23 5.496 0.32 ;
      RECT 5.226 0.78 5.695 0.87 ;
      RECT 5.555 0.759 5.695 0.87 ;
      RECT 2.359 0.17 2.449 0.82 ;
      RECT 5.226 0.456 5.316 0.87 ;
      RECT 4.115 0.456 5.316 0.546 ;
      RECT 4.735 0.266 4.825 0.546 ;
      RECT 4.115 0.17 4.205 0.546 ;
      RECT 3.086 0.265 3.39 0.355 ;
      RECT 3.075 0.221 3.086 0.35 ;
      RECT 3.075 0.265 3.436 0.332 ;
      RECT 3.029 0.193 3.075 0.321 ;
      RECT 3.352 0.246 3.485 0.279 ;
      RECT 3.436 0.175 3.447 0.304 ;
      RECT 2.991 0.246 3.124 0.279 ;
      RECT 3.447 0.17 4.205 0.26 ;
      RECT 2.359 0.17 3.029 0.26 ;
      RECT 3.39 0.204 4.205 0.26 ;
      RECT 3.422 0.96 3.842 1.05 ;
      RECT 3.38 0.901 3.422 1.029 ;
      RECT 3.342 0.96 3.842 0.989 ;
      RECT 2.72 0.88 3.38 0.97 ;
      RECT 2.72 0.941 3.46 0.97 ;
      RECT 2.72 0.739 2.81 0.97 ;
      RECT 3.503 0.7 3.667 0.87 ;
      RECT 3.565 0.36 3.667 0.87 ;
      RECT 2.999 0.7 3.667 0.79 ;
      RECT 3.515 0.36 3.667 0.45 ;
      RECT 2.467 0.959 2.629 1.049 ;
      RECT 2.539 0.35 2.629 1.049 ;
      RECT 3.206 0.52 3.419 0.61 ;
      RECT 2.539 0.445 3.296 0.535 ;
      RECT 2.539 0.35 2.679 0.535 ;
      RECT 1.872 0.96 2.357 1.05 ;
      RECT 1.861 0.916 1.872 1.045 ;
      RECT 0.761 0.935 1.1 1.025 ;
      RECT 1.815 0.888 1.861 1.016 ;
      RECT 2.179 0.208 2.269 1.05 ;
      RECT 1.777 0.941 1.91 0.974 ;
      RECT 1.01 0.865 1.815 0.955 ;
      RECT 1.349 0.325 1.439 0.955 ;
      RECT 1.034 0.325 1.439 0.415 ;
      RECT 1.949 0.78 2.089 0.87 ;
      RECT 1.949 0.27 2.039 0.87 ;
      RECT 1.787 0.27 2.039 0.36 ;
      RECT 0.07 0.201 0.16 1.076 ;
      RECT 0.71 0.445 0.8 0.727 ;
      RECT 0.71 0.561 1.255 0.651 ;
      RECT 0.07 0.445 0.8 0.535 ;
      RECT 4.334 0.661 5.061 0.751 ;
  END
END EDFFQX2H7R

MACRO ESDFFQX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ESDFFQX0P5H7R 0 0 ;
  SIZE 9.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 9.2 1.48 ;
        RECT 8.749 1.095 8.839 1.48 ;
        RECT 8.113 1.095 8.203 1.48 ;
        RECT 7.603 0.987 7.693 1.48 ;
        RECT 5.372 1.24 5.512 1.48 ;
        RECT 4.653 1.24 4.793 1.48 ;
        RECT 3.451 1.24 3.591 1.48 ;
        RECT 1.495 1.07 1.585 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 9.2 0.08 ;
        RECT 8.72 -0.08 8.86 0.36 ;
        RECT 8.199 -0.08 8.289 0.39 ;
        RECT 7.43 -0.08 7.57 0.16 ;
        RECT 5.397 -0.08 5.487 0.301 ;
        RECT 4.57 -0.08 4.71 0.275 ;
        RECT 3.265 -0.08 3.355 0.358 ;
        RECT 1.505 -0.08 1.645 0.305 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 8.65 0.553 8.915 0.808 ;
      LAYER MET2 ;
        RECT 8.65 0.425 8.75 0.96 ;
      LAYER VIA1 ;
        RECT 8.655 0.655 8.745 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.42 0.65 0.575 0.825 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.145 0.45 1.235 0.795 ;
        RECT 0.225 0.45 1.235 0.55 ;
        RECT 0.66 0.45 0.8 0.62 ;
        RECT 0.225 0.45 0.34 0.605 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 8.412 0.245 8.552 0.886 ;
      LAYER MET2 ;
        RECT 8.45 0.23 8.55 0.76 ;
      LAYER VIA1 ;
        RECT 8.455 0.455 8.545 0.545 ;
    END
  END Q
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.825 0.425 2.967 0.58 ;
        RECT 2.265 0.71 2.925 0.8 ;
        RECT 2.825 0.425 2.925 0.8 ;
        RECT 2.265 0.655 2.407 0.8 ;
      LAYER MET2 ;
        RECT 2.85 0.23 2.95 0.76 ;
      LAYER VIA1 ;
        RECT 2.855 0.455 2.945 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.025 0.65 3.285 0.79 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 8.397 1.044 8.571 1.134 ;
      RECT 8.352 0.983 8.397 1.112 ;
      RECT 8.352 1.044 8.617 1.111 ;
      RECT 8.533 1.025 8.662 1.066 ;
      RECT 8.306 1.025 8.435 1.066 ;
      RECT 8.571 0.983 8.662 1.066 ;
      RECT 8.306 0.938 8.352 1.066 ;
      RECT 8.571 0.983 8.7 1.024 ;
      RECT 8.268 0.983 8.397 1.024 ;
      RECT 9.023 0.29 9.113 1.005 ;
      RECT 8.013 0.915 8.306 1.005 ;
      RECT 8.617 0.937 9.113 1.005 ;
      RECT 8.662 0.915 9.113 1.005 ;
      RECT 8.013 0.17 8.103 1.005 ;
      RECT 4.14 0.725 4.33 0.87 ;
      RECT 5.517 0.405 5.607 0.788 ;
      RECT 4.14 0.17 4.23 0.87 ;
      RECT 7.063 0.17 7.153 0.648 ;
      RECT 3.64 0.495 3.755 0.635 ;
      RECT 5.217 0.405 5.667 0.495 ;
      RECT 5.577 0.17 5.667 0.495 ;
      RECT 3.64 0.17 3.73 0.635 ;
      RECT 4.14 0.365 4.897 0.455 ;
      RECT 4.807 0.195 4.897 0.455 ;
      RECT 5.217 0.295 5.307 0.495 ;
      RECT 7.063 0.25 7.648 0.34 ;
      RECT 5.198 0.204 5.217 0.334 ;
      RECT 5.159 0.277 5.298 0.305 ;
      RECT 4.807 0.195 5.198 0.285 ;
      RECT 7.063 0.25 7.728 0.28 ;
      RECT 4.807 0.237 5.263 0.285 ;
      RECT 7.689 0.17 8.103 0.26 ;
      RECT 3.64 0.17 4.23 0.26 ;
      RECT 7.609 0.23 8.103 0.26 ;
      RECT 7.648 0.19 7.689 0.32 ;
      RECT 5.577 0.17 7.153 0.26 ;
      RECT 5.716 1.14 7.513 1.23 ;
      RECT 7.423 0.807 7.513 1.23 ;
      RECT 3.681 1.14 4.532 1.23 ;
      RECT 1.675 1.14 3.332 1.23 ;
      RECT 4.895 1.124 5.244 1.214 ;
      RECT 5.675 1.08 5.716 1.21 ;
      RECT 3.681 1.14 4.573 1.21 ;
      RECT 1.675 1.14 3.373 1.21 ;
      RECT 5.636 1.14 7.513 1.17 ;
      RECT 3.681 1.14 4.612 1.17 ;
      RECT 1.675 1.14 3.412 1.17 ;
      RECT 4.831 1.124 5.308 1.169 ;
      RECT 5.27 1.06 5.675 1.15 ;
      RECT 5.716 1.12 5.755 1.23 ;
      RECT 3.293 1.12 3.771 1.15 ;
      RECT 1.675 0.66 1.765 1.23 ;
      RECT 5.244 1.073 5.27 1.201 ;
      RECT 4.493 1.12 4.933 1.15 ;
      RECT 4.895 1.105 4.933 1.214 ;
      RECT 5.206 1.105 5.716 1.15 ;
      RECT 4.869 1.073 4.895 1.201 ;
      RECT 3.332 1.08 3.771 1.15 ;
      RECT 3.373 1.06 3.771 1.15 ;
      RECT 4.532 1.08 4.895 1.15 ;
      RECT 4.573 1.06 4.869 1.15 ;
      RECT 7.833 0.35 7.923 0.964 ;
      RECT 7.423 0.807 7.923 0.897 ;
      RECT 1.505 0.66 1.765 0.8 ;
      RECT 7.783 0.35 7.923 0.44 ;
      RECT 6.673 0.96 7.333 1.05 ;
      RECT 7.243 0.578 7.333 1.05 ;
      RECT 6.833 0.357 6.923 1.05 ;
      RECT 7.243 0.578 7.648 0.668 ;
      RECT 6.833 0.357 6.973 0.483 ;
      RECT 5.832 0.96 6.563 1.05 ;
      RECT 6.465 0.357 6.563 1.05 ;
      RECT 5.791 0.9 5.832 1.03 ;
      RECT 4.968 0.88 5.127 1.005 ;
      RECT 5.002 0.41 5.127 1.005 ;
      RECT 5.752 0.96 6.563 0.99 ;
      RECT 4.968 0.88 5.791 0.97 ;
      RECT 4.968 0.94 5.871 0.97 ;
      RECT 4.459 0.545 4.574 0.76 ;
      RECT 4.459 0.545 5.127 0.635 ;
      RECT 4.987 0.41 5.127 0.635 ;
      RECT 6.423 0.357 6.563 0.447 ;
      RECT 6.178 0.388 6.318 0.87 ;
      RECT 5.765 0.388 6.318 0.53 ;
      RECT 3.979 0.96 4.448 1.05 ;
      RECT 3.946 0.96 4.448 1.034 ;
      RECT 3.946 0.96 4.489 1.03 ;
      RECT 3.9 0.96 4.489 0.994 ;
      RECT 3.9 0.96 4.528 0.99 ;
      RECT 3.899 0.35 3.989 0.971 ;
      RECT 4.664 0.725 4.754 0.97 ;
      RECT 4.409 0.94 4.754 0.97 ;
      RECT 4.489 0.88 4.754 0.97 ;
      RECT 3.899 0.945 4.018 0.971 ;
      RECT 4.448 0.9 4.754 0.97 ;
      RECT 4.664 0.725 4.893 0.815 ;
      RECT 3.84 0.35 3.989 0.44 ;
      RECT 2.53 0.901 3.313 0.991 ;
      RECT 2.53 0.901 3.334 0.981 ;
      RECT 3.375 0.448 3.465 0.97 ;
      RECT 3.275 0.89 3.465 0.97 ;
      RECT 3.296 0.88 3.465 0.97 ;
      RECT 3.085 0.448 3.465 0.538 ;
      RECT 3.085 0.233 3.175 0.538 ;
      RECT 2.68 0.216 3.14 0.306 ;
      RECT 2.035 0.78 2.175 0.87 ;
      RECT 2.035 0.357 2.125 0.87 ;
      RECT 2.58 0.418 2.72 0.62 ;
      RECT 2.035 0.418 2.72 0.508 ;
      RECT 2.035 0.357 2.175 0.508 ;
      RECT 1.01 1.095 1.229 1.185 ;
      RECT 1.139 0.915 1.229 1.185 ;
      RECT 1.855 0.96 2.42 1.05 ;
      RECT 1.139 0.915 1.289 1.005 ;
      RECT 1.855 0.17 1.945 1.05 ;
      RECT 1.251 0.896 1.371 0.946 ;
      RECT 1.289 0.859 1.325 0.987 ;
      RECT 1.325 0.267 1.415 0.901 ;
      RECT 1.325 0.395 1.945 0.485 ;
      RECT 1.835 0.17 1.945 0.485 ;
      RECT 0.76 0.267 1.415 0.357 ;
      RECT 2.295 0.17 2.435 0.306 ;
      RECT 1.835 0.17 2.435 0.26 ;
      RECT 0.045 0.915 0.181 1.121 ;
      RECT 0.045 0.915 1.005 1.005 ;
      RECT 0.915 0.655 1.005 1.005 ;
      RECT 0.045 0.232 0.135 1.121 ;
      RECT 0.045 0.232 0.16 0.372 ;
  END
END ESDFFQX0P5H7R

MACRO ESDFFQX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ESDFFQX1H7R 0 0 ;
  SIZE 9.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 9.2 1.48 ;
        RECT 8.749 1.095 8.839 1.48 ;
        RECT 8.113 1.095 8.203 1.48 ;
        RECT 7.603 0.987 7.693 1.48 ;
        RECT 5.278 1.24 5.418 1.48 ;
        RECT 4.653 1.24 4.793 1.48 ;
        RECT 3.451 1.24 3.591 1.48 ;
        RECT 1.495 1.07 1.585 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 9.2 0.08 ;
        RECT 8.72 -0.08 8.86 0.36 ;
        RECT 8.199 -0.08 8.289 0.39 ;
        RECT 7.43 -0.08 7.57 0.16 ;
        RECT 5.397 -0.08 5.487 0.301 ;
        RECT 4.57 -0.08 4.71 0.275 ;
        RECT 3.265 -0.08 3.355 0.358 ;
        RECT 1.505 -0.08 1.645 0.305 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 8.65 0.553 8.915 0.808 ;
      LAYER MET2 ;
        RECT 8.65 0.425 8.75 0.96 ;
      LAYER VIA1 ;
        RECT 8.655 0.655 8.745 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.65 0.575 0.75 ;
        RECT 0.36 0.695 0.551 0.814 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.145 0.465 1.235 0.795 ;
        RECT 0.225 0.465 1.235 0.555 ;
        RECT 0.66 0.465 0.8 0.62 ;
        RECT 0.225 0.45 0.375 0.555 ;
        RECT 0.225 0.45 0.34 0.605 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 8.412 0.245 8.552 0.886 ;
      LAYER MET2 ;
        RECT 8.45 0.23 8.55 0.76 ;
      LAYER VIA1 ;
        RECT 8.455 0.455 8.545 0.545 ;
    END
  END Q
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.825 0.425 2.967 0.58 ;
        RECT 2.265 0.71 2.925 0.8 ;
        RECT 2.825 0.425 2.925 0.8 ;
        RECT 2.265 0.655 2.407 0.8 ;
      LAYER MET2 ;
        RECT 2.85 0.23 2.95 0.76 ;
      LAYER VIA1 ;
        RECT 2.855 0.455 2.945 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.025 0.65 3.285 0.79 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 8.397 1.044 8.571 1.134 ;
      RECT 8.352 0.983 8.397 1.112 ;
      RECT 8.352 1.044 8.617 1.111 ;
      RECT 8.533 1.025 8.662 1.066 ;
      RECT 8.306 1.025 8.435 1.066 ;
      RECT 8.571 0.983 8.662 1.066 ;
      RECT 8.306 0.938 8.352 1.066 ;
      RECT 8.571 0.983 8.7 1.024 ;
      RECT 8.268 0.983 8.397 1.024 ;
      RECT 9.023 0.29 9.113 1.005 ;
      RECT 8.013 0.915 8.306 1.005 ;
      RECT 8.617 0.937 9.113 1.005 ;
      RECT 8.662 0.915 9.113 1.005 ;
      RECT 8.013 0.17 8.103 1.005 ;
      RECT 4.14 0.725 4.33 0.87 ;
      RECT 5.517 0.405 5.607 0.788 ;
      RECT 4.14 0.17 4.23 0.87 ;
      RECT 7.063 0.17 7.153 0.648 ;
      RECT 3.64 0.495 3.755 0.635 ;
      RECT 5.217 0.405 5.667 0.495 ;
      RECT 5.577 0.17 5.667 0.495 ;
      RECT 3.64 0.17 3.73 0.635 ;
      RECT 4.14 0.365 4.897 0.455 ;
      RECT 4.807 0.195 4.897 0.455 ;
      RECT 5.217 0.295 5.307 0.495 ;
      RECT 7.063 0.25 7.648 0.34 ;
      RECT 5.198 0.204 5.217 0.334 ;
      RECT 5.159 0.277 5.298 0.305 ;
      RECT 4.807 0.195 5.198 0.285 ;
      RECT 7.063 0.25 7.728 0.28 ;
      RECT 4.807 0.237 5.263 0.285 ;
      RECT 7.689 0.17 8.103 0.26 ;
      RECT 3.64 0.17 4.23 0.26 ;
      RECT 7.609 0.23 8.103 0.26 ;
      RECT 7.648 0.19 7.689 0.32 ;
      RECT 5.577 0.17 7.153 0.26 ;
      RECT 5.716 1.14 7.513 1.23 ;
      RECT 7.423 0.807 7.513 1.23 ;
      RECT 3.681 1.14 4.532 1.23 ;
      RECT 1.675 1.14 3.332 1.23 ;
      RECT 5.675 1.14 7.513 1.21 ;
      RECT 3.681 1.14 4.573 1.21 ;
      RECT 1.675 1.14 3.373 1.21 ;
      RECT 5.636 1.14 7.513 1.17 ;
      RECT 3.681 1.14 4.612 1.17 ;
      RECT 1.675 1.14 3.412 1.17 ;
      RECT 4.573 1.06 5.675 1.15 ;
      RECT 4.493 1.12 5.755 1.15 ;
      RECT 3.293 1.12 3.771 1.15 ;
      RECT 1.675 0.66 1.765 1.23 ;
      RECT 4.532 1.08 5.716 1.15 ;
      RECT 3.332 1.08 3.771 1.15 ;
      RECT 3.373 1.06 3.771 1.15 ;
      RECT 7.833 0.35 7.923 0.964 ;
      RECT 7.423 0.807 7.923 0.897 ;
      RECT 1.505 0.66 1.765 0.8 ;
      RECT 7.783 0.35 7.923 0.44 ;
      RECT 6.673 0.96 7.333 1.05 ;
      RECT 7.243 0.578 7.333 1.05 ;
      RECT 6.833 0.357 6.923 1.05 ;
      RECT 7.243 0.578 7.648 0.668 ;
      RECT 6.833 0.357 6.973 0.483 ;
      RECT 5.832 0.96 6.563 1.05 ;
      RECT 6.465 0.357 6.563 1.05 ;
      RECT 5.791 0.9 5.832 1.03 ;
      RECT 5.752 0.96 6.563 0.99 ;
      RECT 4.968 0.88 5.791 0.97 ;
      RECT 4.968 0.94 5.871 0.97 ;
      RECT 5.002 0.398 5.127 0.97 ;
      RECT 4.459 0.545 4.574 0.76 ;
      RECT 4.459 0.545 5.127 0.635 ;
      RECT 4.987 0.398 5.127 0.635 ;
      RECT 6.423 0.357 6.563 0.447 ;
      RECT 6.178 0.388 6.318 0.87 ;
      RECT 5.765 0.388 6.318 0.53 ;
      RECT 3.979 0.96 4.448 1.05 ;
      RECT 3.946 0.96 4.448 1.034 ;
      RECT 3.946 0.96 4.489 1.03 ;
      RECT 3.9 0.96 4.489 0.994 ;
      RECT 3.9 0.96 4.528 0.99 ;
      RECT 3.899 0.35 3.989 0.971 ;
      RECT 4.664 0.725 4.754 0.97 ;
      RECT 4.409 0.94 4.754 0.97 ;
      RECT 4.489 0.88 4.754 0.97 ;
      RECT 3.899 0.945 4.018 0.971 ;
      RECT 4.448 0.9 4.754 0.97 ;
      RECT 4.664 0.725 4.893 0.815 ;
      RECT 3.84 0.35 3.989 0.44 ;
      RECT 2.53 0.901 3.313 0.991 ;
      RECT 2.53 0.901 3.334 0.981 ;
      RECT 3.375 0.448 3.465 0.97 ;
      RECT 3.275 0.89 3.465 0.97 ;
      RECT 3.296 0.88 3.465 0.97 ;
      RECT 3.085 0.448 3.465 0.538 ;
      RECT 3.085 0.233 3.175 0.538 ;
      RECT 2.68 0.216 3.14 0.306 ;
      RECT 2.035 0.78 2.175 0.87 ;
      RECT 2.035 0.357 2.125 0.87 ;
      RECT 2.58 0.418 2.72 0.62 ;
      RECT 2.035 0.418 2.72 0.508 ;
      RECT 2.035 0.357 2.175 0.508 ;
      RECT 1.01 1.095 1.229 1.185 ;
      RECT 1.139 0.915 1.229 1.185 ;
      RECT 1.855 0.96 2.42 1.05 ;
      RECT 1.139 0.915 1.289 1.005 ;
      RECT 1.855 0.17 1.945 1.05 ;
      RECT 1.251 0.896 1.371 0.946 ;
      RECT 1.289 0.859 1.325 0.987 ;
      RECT 1.325 0.267 1.415 0.901 ;
      RECT 1.325 0.395 1.945 0.485 ;
      RECT 1.835 0.17 1.945 0.485 ;
      RECT 0.76 0.267 1.415 0.357 ;
      RECT 2.295 0.17 2.435 0.306 ;
      RECT 1.835 0.17 2.435 0.26 ;
      RECT 0.045 0.915 0.181 1.121 ;
      RECT 0.045 0.915 1.005 1.005 ;
      RECT 0.915 0.655 1.005 1.005 ;
      RECT 0.045 0.232 0.135 1.121 ;
      RECT 0.045 0.232 0.16 0.372 ;
  END
END ESDFFQX1H7R

MACRO ESDFFQX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ESDFFQX2H7R 0 0 ;
  SIZE 9.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 9.2 1.48 ;
        RECT 8.749 1.095 8.839 1.48 ;
        RECT 8.113 1.095 8.203 1.48 ;
        RECT 7.603 0.987 7.693 1.48 ;
        RECT 5.278 1.24 5.418 1.48 ;
        RECT 4.653 1.24 4.793 1.48 ;
        RECT 3.451 1.24 3.591 1.48 ;
        RECT 1.495 1.07 1.585 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 9.2 0.08 ;
        RECT 8.72 -0.08 8.86 0.365 ;
        RECT 8.199 -0.08 8.289 0.39 ;
        RECT 7.43 -0.08 7.57 0.16 ;
        RECT 5.397 -0.08 5.487 0.301 ;
        RECT 4.57 -0.08 4.71 0.275 ;
        RECT 3.24 -0.08 3.38 0.333 ;
        RECT 1.505 -0.08 1.645 0.305 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 8.65 0.553 8.915 0.808 ;
      LAYER MET2 ;
        RECT 8.65 0.425 8.75 0.96 ;
      LAYER VIA1 ;
        RECT 8.655 0.655 8.745 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.36 0.695 0.575 0.814 ;
        RECT 0.425 0.65 0.575 0.814 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.145 0.45 1.235 0.795 ;
        RECT 0.225 0.45 1.235 0.555 ;
        RECT 0.66 0.45 0.8 0.62 ;
        RECT 0.225 0.45 0.34 0.605 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 8.412 0.25 8.552 0.886 ;
      LAYER MET2 ;
        RECT 8.45 0.23 8.55 0.76 ;
      LAYER VIA1 ;
        RECT 8.455 0.455 8.545 0.545 ;
    END
  END Q
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.825 0.425 2.967 0.58 ;
        RECT 2.265 0.71 2.925 0.8 ;
        RECT 2.825 0.425 2.925 0.8 ;
        RECT 2.265 0.655 2.407 0.8 ;
      LAYER MET2 ;
        RECT 2.85 0.23 2.95 0.76 ;
      LAYER VIA1 ;
        RECT 2.855 0.455 2.945 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.05 0.625 3.285 0.79 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 8.397 1.044 8.571 1.134 ;
      RECT 8.352 0.983 8.397 1.112 ;
      RECT 8.352 1.044 8.617 1.111 ;
      RECT 8.533 1.025 8.662 1.066 ;
      RECT 8.306 1.025 8.435 1.066 ;
      RECT 8.571 0.983 8.662 1.066 ;
      RECT 8.306 0.938 8.352 1.066 ;
      RECT 8.571 0.983 8.7 1.024 ;
      RECT 8.268 0.983 8.397 1.024 ;
      RECT 9.023 0.29 9.113 1.005 ;
      RECT 8.013 0.915 8.306 1.005 ;
      RECT 8.617 0.937 9.113 1.005 ;
      RECT 8.662 0.915 9.113 1.005 ;
      RECT 8.013 0.17 8.103 1.005 ;
      RECT 4.14 0.725 4.33 0.87 ;
      RECT 5.517 0.405 5.607 0.788 ;
      RECT 4.14 0.17 4.23 0.87 ;
      RECT 7.063 0.17 7.153 0.648 ;
      RECT 3.64 0.495 3.755 0.635 ;
      RECT 5.217 0.405 5.667 0.495 ;
      RECT 5.577 0.17 5.667 0.495 ;
      RECT 3.64 0.17 3.73 0.635 ;
      RECT 4.14 0.365 4.897 0.455 ;
      RECT 4.807 0.195 4.897 0.455 ;
      RECT 5.217 0.295 5.307 0.495 ;
      RECT 7.063 0.25 7.648 0.34 ;
      RECT 5.198 0.204 5.217 0.334 ;
      RECT 5.159 0.277 5.298 0.305 ;
      RECT 4.807 0.195 5.198 0.285 ;
      RECT 7.063 0.25 7.728 0.28 ;
      RECT 4.807 0.237 5.263 0.285 ;
      RECT 7.689 0.17 8.103 0.26 ;
      RECT 3.64 0.17 4.23 0.26 ;
      RECT 7.609 0.23 8.103 0.26 ;
      RECT 7.648 0.19 7.689 0.32 ;
      RECT 5.577 0.17 7.153 0.26 ;
      RECT 5.716 1.14 7.513 1.23 ;
      RECT 7.423 0.807 7.513 1.23 ;
      RECT 3.681 1.14 4.532 1.23 ;
      RECT 1.675 1.14 3.332 1.23 ;
      RECT 5.675 1.14 7.513 1.21 ;
      RECT 3.681 1.14 4.573 1.21 ;
      RECT 1.675 1.14 3.373 1.21 ;
      RECT 5.636 1.14 7.513 1.17 ;
      RECT 3.681 1.14 4.612 1.17 ;
      RECT 1.675 1.14 3.412 1.17 ;
      RECT 4.573 1.06 5.675 1.15 ;
      RECT 4.493 1.12 5.755 1.15 ;
      RECT 3.293 1.12 3.771 1.15 ;
      RECT 1.675 0.66 1.765 1.23 ;
      RECT 4.532 1.08 5.716 1.15 ;
      RECT 3.332 1.08 3.771 1.15 ;
      RECT 3.373 1.06 3.771 1.15 ;
      RECT 7.833 0.35 7.923 0.964 ;
      RECT 7.423 0.807 7.923 0.897 ;
      RECT 1.505 0.66 1.765 0.8 ;
      RECT 7.783 0.35 7.923 0.44 ;
      RECT 6.673 0.96 7.333 1.05 ;
      RECT 7.243 0.578 7.333 1.05 ;
      RECT 6.833 0.357 6.923 1.05 ;
      RECT 7.243 0.578 7.648 0.668 ;
      RECT 6.833 0.357 6.973 0.483 ;
      RECT 5.832 0.96 6.563 1.05 ;
      RECT 6.465 0.357 6.563 1.05 ;
      RECT 5.791 0.9 5.832 1.03 ;
      RECT 5.752 0.96 6.563 0.99 ;
      RECT 4.968 0.88 5.791 0.97 ;
      RECT 4.968 0.94 5.871 0.97 ;
      RECT 5.002 0.398 5.127 0.97 ;
      RECT 4.459 0.545 4.574 0.76 ;
      RECT 4.459 0.545 5.127 0.635 ;
      RECT 4.987 0.398 5.127 0.635 ;
      RECT 6.423 0.357 6.563 0.447 ;
      RECT 6.178 0.388 6.318 0.87 ;
      RECT 5.765 0.388 6.318 0.53 ;
      RECT 3.979 0.96 4.448 1.05 ;
      RECT 3.946 0.96 4.448 1.034 ;
      RECT 3.946 0.96 4.489 1.03 ;
      RECT 3.9 0.96 4.489 0.994 ;
      RECT 3.9 0.96 4.528 0.99 ;
      RECT 3.899 0.35 3.989 0.971 ;
      RECT 4.664 0.725 4.754 0.97 ;
      RECT 4.409 0.94 4.754 0.97 ;
      RECT 4.489 0.88 4.754 0.97 ;
      RECT 3.899 0.945 4.018 0.971 ;
      RECT 4.448 0.9 4.754 0.97 ;
      RECT 4.664 0.725 4.893 0.815 ;
      RECT 3.84 0.35 3.989 0.44 ;
      RECT 2.53 0.901 3.313 0.991 ;
      RECT 2.53 0.901 3.334 0.981 ;
      RECT 3.375 0.445 3.465 0.97 ;
      RECT 3.275 0.89 3.465 0.97 ;
      RECT 3.296 0.88 3.465 0.97 ;
      RECT 3.06 0.445 3.465 0.535 ;
      RECT 3.06 0.221 3.15 0.535 ;
      RECT 2.68 0.216 3.14 0.306 ;
      RECT 2.035 0.78 2.175 0.87 ;
      RECT 2.035 0.357 2.125 0.87 ;
      RECT 2.58 0.418 2.72 0.62 ;
      RECT 2.035 0.418 2.72 0.508 ;
      RECT 2.035 0.357 2.175 0.508 ;
      RECT 1.01 1.095 1.229 1.185 ;
      RECT 1.139 0.915 1.229 1.185 ;
      RECT 1.855 0.96 2.42 1.05 ;
      RECT 1.139 0.915 1.289 1.005 ;
      RECT 1.855 0.17 1.945 1.05 ;
      RECT 1.251 0.896 1.371 0.946 ;
      RECT 1.289 0.859 1.325 0.987 ;
      RECT 1.325 0.267 1.415 0.901 ;
      RECT 1.325 0.395 1.945 0.485 ;
      RECT 0.76 0.267 1.415 0.357 ;
      RECT 2.295 0.17 2.435 0.306 ;
      RECT 1.855 0.17 2.435 0.26 ;
      RECT 0.045 0.915 0.181 1.121 ;
      RECT 0.045 0.915 1.005 1.005 ;
      RECT 0.915 0.655 1.005 1.005 ;
      RECT 0.045 0.232 0.135 1.121 ;
      RECT 0.045 0.232 0.16 0.372 ;
  END
END ESDFFQX2H7R

MACRO FILLCAP16H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILLCAP16H7R 0 0 ;
  SIZE 3.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.2 1.48 ;
        RECT 0.07 1.045 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.2 0.08 ;
        RECT 3.04 -0.08 3.13 0.355 ;
    END
  END VSS
  OBS
    LAYER MET1 ;
      RECT 3.04 0.445 3.13 1.045 ;
      RECT 0.25 0.445 3.13 0.58 ;
      RECT 0.07 0.72 2.94 0.86 ;
      RECT 0.07 0.255 0.16 0.86 ;
  END
END FILLCAP16H7R

MACRO FILLCAP32H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILLCAP32H7R 0 0 ;
  SIZE 6.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.4 1.48 ;
        RECT 0.07 1.045 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.4 0.08 ;
        RECT 6.24 -0.08 6.33 0.355 ;
    END
  END VSS
  OBS
    LAYER MET1 ;
      RECT 6.24 0.445 6.33 1.045 ;
      RECT 0.25 0.445 6.33 0.585 ;
      RECT 0.07 0.72 6.14 0.86 ;
      RECT 0.07 0.255 0.16 0.86 ;
  END
END FILLCAP32H7R

MACRO FILLCAP4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILLCAP4H7R 0 0 ;
  SIZE 0.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.8 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.8 0.08 ;
        RECT 0.64 -0.08 0.73 0.345 ;
    END
  END VSS
  OBS
    LAYER MET1 ;
      RECT 0.64 0.465 0.73 1.045 ;
      RECT 0.25 0.465 0.73 0.605 ;
      RECT 0.07 0.72 0.54 0.86 ;
      RECT 0.07 0.255 0.16 0.86 ;
  END
END FILLCAP4H7R

MACRO FILLCAP8H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILLCAP8H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.07 1.045 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.44 -0.08 1.53 0.355 ;
    END
  END VSS
  OBS
    LAYER MET1 ;
      RECT 1.44 0.445 1.53 1.045 ;
      RECT 0.25 0.445 1.53 0.58 ;
      RECT 0.07 0.72 1.34 0.86 ;
      RECT 0.07 0.255 0.16 0.86 ;
  END
END FILLCAP8H7R

MACRO FILLER16H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILLER16H7R 0 0 ;
  SIZE 3.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.2 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.2 0.08 ;
    END
  END VSS
END FILLER16H7R

MACRO FILLER1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILLER1H7R 0 0 ;
  SIZE 0.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.2 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.2 0.08 ;
    END
  END VSS
END FILLER1H7R

MACRO FILLER2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILLER2H7R 0 0 ;
  SIZE 0.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.4 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.4 0.08 ;
    END
  END VSS
END FILLER2H7R

MACRO FILLER32H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILLER32H7R 0 0 ;
  SIZE 6.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.4 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.4 0.08 ;
    END
  END VSS
END FILLER32H7R

MACRO FILLER4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILLER4H7R 0 0 ;
  SIZE 0.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.8 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.8 0.08 ;
    END
  END VSS
END FILLER4H7R

MACRO FILLER64H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILLER64H7R 0 0 ;
  SIZE 12.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 12.8 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 12.8 0.08 ;
    END
  END VSS
END FILLER64H7R

MACRO FILLER8H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILLER8H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
    END
  END VSS
END FILLER8H7R

MACRO FILLTAPH7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILLTAPH7R 0 0 ;
  SIZE 0.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.4 1.48 ;
        RECT 0.055 0.66 0.345 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.4 0.08 ;
        RECT 0.055 -0.08 0.345 0.57 ;
    END
  END VSS
END FILLTAPH7R

MACRO ICGNX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGNX0P5H7R 0 0 ;
  SIZE 4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4 1.48 ;
        RECT 3.275 1.075 3.415 1.48 ;
        RECT 2.245 1.24 2.385 1.48 ;
        RECT 1.495 1.095 1.635 1.48 ;
        RECT 0.32 1.05 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4 0.08 ;
        RECT 3.31 -0.08 3.45 0.305 ;
        RECT 2.55 -0.08 2.69 0.16 ;
        RECT 1.556 -0.08 1.696 0.16 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 2.45 0.51 2.79 0.6 ;
        RECT 2.625 0.455 2.79 0.6 ;
      LAYER MET2 ;
        RECT 2.65 0.23 2.75 0.76 ;
      LAYER VIA1 ;
        RECT 2.655 0.455 2.745 0.545 ;
    END
  END CKN
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.395 0.625 1.545 0.805 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END E
  PIN ECK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.54 1.075 3.916 1.165 ;
        RECT 3.826 0.255 3.916 1.165 ;
        RECT 3.56 0.255 3.916 0.345 ;
      LAYER MET2 ;
        RECT 3.65 0.18 3.75 0.56 ;
      LAYER VIA1 ;
        RECT 3.655 0.255 3.745 0.345 ;
    END
  END ECK
  OBS
    LAYER MET1 ;
      RECT 2.503 1.14 3.125 1.23 ;
      RECT 3.035 0.89 3.125 1.23 ;
      RECT 2.497 1.099 2.503 1.227 ;
      RECT 2.451 1.073 2.497 1.201 ;
      RECT 0.68 1.1 1.23 1.19 ;
      RECT 1.14 0.53 1.23 1.19 ;
      RECT 2.413 1.14 3.125 1.159 ;
      RECT 1.725 1.05 2.451 1.14 ;
      RECT 1.725 1.121 2.541 1.14 ;
      RECT 0.68 0.825 0.77 1.19 ;
      RECT 1.725 0.915 1.815 1.14 ;
      RECT 1.14 0.915 1.815 1.005 ;
      RECT 3.035 0.89 3.736 0.98 ;
      RECT 3.646 0.48 3.736 0.98 ;
      RECT 1.14 0.53 1.286 0.62 ;
      RECT 3.293 0.48 3.736 0.57 ;
      RECT 3.267 0.429 3.293 0.557 ;
      RECT 3.221 0.393 3.267 0.521 ;
      RECT 3.221 0.461 3.331 0.521 ;
      RECT 3.175 0.347 3.221 0.475 ;
      RECT 3.131 0.205 3.175 0.43 ;
      RECT 3.085 0.205 3.175 0.385 ;
      RECT 1.985 0.87 2.305 0.96 ;
      RECT 2.215 0.35 2.305 0.96 ;
      RECT 2.215 0.71 3.556 0.8 ;
      RECT 3.466 0.66 3.556 0.8 ;
      RECT 2.215 0.35 2.355 0.44 ;
      RECT 1.675 0.69 2.125 0.78 ;
      RECT 2.035 0.17 2.125 0.78 ;
      RECT 1.675 0.43 1.765 0.78 ;
      RECT 2.9 0.485 3.08 0.575 ;
      RECT 0.76 0.445 0.941 0.535 ;
      RECT 1.404 0.43 1.765 0.52 ;
      RECT 1.362 0.371 1.404 0.499 ;
      RECT 2.9 0.25 2.99 0.575 ;
      RECT 1.324 0.43 1.765 0.459 ;
      RECT 0.903 0.426 1.036 0.459 ;
      RECT 0.987 0.355 0.998 0.484 ;
      RECT 0.998 0.35 1.362 0.44 ;
      RECT 1.404 0.411 1.442 0.52 ;
      RECT 0.941 0.384 0.987 0.512 ;
      RECT 2.473 0.25 2.99 0.34 ;
      RECT 2.431 0.191 2.473 0.319 ;
      RECT 2.393 0.25 2.99 0.279 ;
      RECT 2.035 0.17 2.431 0.26 ;
      RECT 2.035 0.231 2.511 0.26 ;
      RECT 0.91 0.645 1 1.01 ;
      RECT 0.225 0.77 0.492 0.86 ;
      RECT 0.225 0.77 0.538 0.837 ;
      RECT 0.454 0.751 0.58 0.793 ;
      RECT 0.225 0.715 0.315 0.86 ;
      RECT 0.492 0.709 0.617 0.754 ;
      RECT 0.538 0.665 0.58 0.793 ;
      RECT 0.58 0.645 1 0.735 ;
      RECT 0.58 0.215 0.67 0.735 ;
      RECT 1.855 0.25 1.945 0.6 ;
      RECT 1.48 0.25 1.945 0.34 ;
      RECT 1.438 0.191 1.48 0.319 ;
      RECT 0.58 0.215 0.915 0.305 ;
      RECT 1.4 0.25 1.945 0.279 ;
      RECT 0.825 0.17 1.438 0.26 ;
      RECT 0.58 0.231 1.518 0.26 ;
      RECT 0.045 0.945 0.185 1.035 ;
      RECT 0.045 0.28 0.135 1.035 ;
      RECT 0.4 0.465 0.49 0.605 ;
      RECT 0.045 0.465 0.49 0.555 ;
      RECT 0.045 0.28 0.185 0.37 ;
      RECT 2.55 0.89 2.92 1.02 ;
  END
END ICGNX0P5H7R

MACRO ICGNX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGNX1H7R 0 0 ;
  SIZE 4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4 1.48 ;
        RECT 3.275 1.075 3.415 1.48 ;
        RECT 2.245 1.24 2.385 1.48 ;
        RECT 1.495 1.095 1.635 1.48 ;
        RECT 0.32 1.05 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4 0.08 ;
        RECT 3.31 -0.08 3.45 0.305 ;
        RECT 2.55 -0.08 2.69 0.16 ;
        RECT 1.556 -0.08 1.696 0.16 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 2.45 0.51 2.79 0.6 ;
        RECT 2.625 0.455 2.79 0.6 ;
      LAYER MET2 ;
        RECT 2.65 0.23 2.75 0.76 ;
      LAYER VIA1 ;
        RECT 2.655 0.455 2.745 0.545 ;
    END
  END CKN
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.395 0.625 1.545 0.805 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END E
  PIN ECK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.54 1.075 3.916 1.165 ;
        RECT 3.826 0.255 3.916 1.165 ;
        RECT 3.56 0.255 3.916 0.345 ;
      LAYER MET2 ;
        RECT 3.65 0.18 3.75 0.56 ;
      LAYER VIA1 ;
        RECT 3.655 0.255 3.745 0.345 ;
    END
  END ECK
  OBS
    LAYER MET1 ;
      RECT 2.503 1.14 3.125 1.23 ;
      RECT 3.035 0.89 3.125 1.23 ;
      RECT 2.497 1.099 2.503 1.227 ;
      RECT 2.451 1.073 2.497 1.201 ;
      RECT 0.68 1.1 1.23 1.19 ;
      RECT 1.14 0.53 1.23 1.19 ;
      RECT 2.413 1.14 3.125 1.159 ;
      RECT 1.725 1.05 2.451 1.14 ;
      RECT 1.725 1.121 2.541 1.14 ;
      RECT 0.68 0.825 0.77 1.19 ;
      RECT 1.725 0.915 1.815 1.14 ;
      RECT 1.14 0.915 1.815 1.005 ;
      RECT 3.035 0.89 3.736 0.98 ;
      RECT 3.646 0.48 3.736 0.98 ;
      RECT 1.14 0.53 1.286 0.62 ;
      RECT 3.293 0.48 3.736 0.57 ;
      RECT 3.267 0.429 3.293 0.557 ;
      RECT 3.221 0.393 3.267 0.521 ;
      RECT 3.221 0.461 3.331 0.521 ;
      RECT 3.175 0.347 3.221 0.475 ;
      RECT 3.131 0.205 3.175 0.43 ;
      RECT 3.085 0.205 3.175 0.385 ;
      RECT 1.955 0.87 2.305 0.96 ;
      RECT 2.215 0.35 2.305 0.96 ;
      RECT 2.215 0.71 3.556 0.8 ;
      RECT 3.466 0.66 3.556 0.8 ;
      RECT 2.215 0.35 2.355 0.44 ;
      RECT 1.675 0.69 2.125 0.78 ;
      RECT 2.035 0.17 2.125 0.78 ;
      RECT 1.675 0.43 1.765 0.78 ;
      RECT 2.9 0.485 3.08 0.575 ;
      RECT 0.76 0.445 0.941 0.535 ;
      RECT 1.404 0.43 1.765 0.52 ;
      RECT 1.362 0.371 1.404 0.499 ;
      RECT 2.9 0.25 2.99 0.575 ;
      RECT 1.324 0.43 1.765 0.459 ;
      RECT 0.903 0.426 1.036 0.459 ;
      RECT 0.987 0.355 0.998 0.484 ;
      RECT 0.998 0.35 1.362 0.44 ;
      RECT 1.404 0.411 1.442 0.52 ;
      RECT 0.941 0.384 0.987 0.512 ;
      RECT 2.473 0.25 2.99 0.34 ;
      RECT 2.431 0.191 2.473 0.319 ;
      RECT 2.393 0.25 2.99 0.279 ;
      RECT 2.035 0.17 2.431 0.26 ;
      RECT 2.035 0.231 2.511 0.26 ;
      RECT 0.91 0.645 1 1.01 ;
      RECT 0.225 0.77 0.492 0.86 ;
      RECT 0.225 0.77 0.538 0.837 ;
      RECT 0.454 0.751 0.58 0.793 ;
      RECT 0.225 0.715 0.315 0.86 ;
      RECT 0.492 0.709 0.617 0.754 ;
      RECT 0.538 0.665 0.58 0.793 ;
      RECT 0.58 0.645 1 0.735 ;
      RECT 0.58 0.215 0.67 0.735 ;
      RECT 1.855 0.25 1.945 0.6 ;
      RECT 1.48 0.25 1.945 0.34 ;
      RECT 1.438 0.191 1.48 0.319 ;
      RECT 0.58 0.215 0.915 0.305 ;
      RECT 1.4 0.25 1.945 0.279 ;
      RECT 0.825 0.17 1.438 0.26 ;
      RECT 0.58 0.231 1.518 0.26 ;
      RECT 0.045 0.945 0.185 1.035 ;
      RECT 0.045 0.275 0.135 1.035 ;
      RECT 0.4 0.465 0.49 0.605 ;
      RECT 0.045 0.465 0.49 0.555 ;
      RECT 0.045 0.275 0.185 0.365 ;
      RECT 2.55 0.93 2.92 1.02 ;
  END
END ICGNX1H7R

MACRO ICGNX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGNX2H7R 0 0 ;
  SIZE 4.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.2 1.48 ;
        RECT 3.88 1.24 4.02 1.48 ;
        RECT 3.275 1.07 3.415 1.48 ;
        RECT 2.245 1.24 2.385 1.48 ;
        RECT 1.495 1.095 1.635 1.48 ;
        RECT 0.32 1.05 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.2 0.08 ;
        RECT 3.825 -0.08 3.965 0.235 ;
        RECT 3.31 -0.08 3.45 0.365 ;
        RECT 2.55 -0.08 2.69 0.16 ;
        RECT 1.556 -0.08 1.696 0.16 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 2.45 0.51 2.79 0.6 ;
        RECT 2.625 0.455 2.79 0.6 ;
      LAYER MET2 ;
        RECT 2.65 0.23 2.75 0.76 ;
      LAYER VIA1 ;
        RECT 2.655 0.455 2.745 0.545 ;
    END
  END CKN
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.41 0.625 1.545 0.825 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END E
  PIN ECK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.855 0.325 3.945 1.069 ;
        RECT 3.54 1.065 3.901 1.114 ;
        RECT 3.799 1.046 3.945 1.069 ;
        RECT 3.837 1.018 3.855 1.146 ;
        RECT 3.585 0.325 3.945 0.415 ;
        RECT 3.54 1.065 3.837 1.155 ;
        RECT 3.585 0.255 3.675 0.415 ;
      LAYER MET2 ;
        RECT 3.85 0.23 3.95 0.76 ;
      LAYER VIA1 ;
        RECT 3.855 0.455 3.945 0.545 ;
    END
  END ECK
  OBS
    LAYER MET1 ;
      RECT 2.503 1.14 3.125 1.23 ;
      RECT 3.035 0.885 3.125 1.23 ;
      RECT 2.497 1.099 2.503 1.227 ;
      RECT 2.451 1.073 2.497 1.201 ;
      RECT 0.68 1.1 1.23 1.19 ;
      RECT 1.14 0.53 1.23 1.19 ;
      RECT 2.413 1.14 3.125 1.159 ;
      RECT 1.725 1.05 2.451 1.14 ;
      RECT 1.725 1.121 2.541 1.14 ;
      RECT 0.68 0.825 0.77 1.19 ;
      RECT 1.725 0.915 1.815 1.14 ;
      RECT 1.14 0.915 1.815 1.005 ;
      RECT 3.035 0.885 3.761 0.975 ;
      RECT 3.671 0.505 3.761 0.975 ;
      RECT 1.14 0.53 1.286 0.62 ;
      RECT 3.278 0.505 3.761 0.595 ;
      RECT 3.267 0.461 3.278 0.59 ;
      RECT 3.221 0.433 3.267 0.561 ;
      RECT 3.175 0.387 3.221 0.515 ;
      RECT 3.175 0.486 3.316 0.515 ;
      RECT 3.131 0.205 3.175 0.47 ;
      RECT 3.085 0.205 3.175 0.425 ;
      RECT 1.985 0.87 2.305 0.96 ;
      RECT 2.215 0.35 2.305 0.96 ;
      RECT 2.215 0.705 3.581 0.795 ;
      RECT 2.215 0.35 2.355 0.44 ;
      RECT 1.675 0.69 2.125 0.78 ;
      RECT 2.035 0.17 2.125 0.78 ;
      RECT 1.675 0.43 1.765 0.78 ;
      RECT 2.9 0.525 3.08 0.615 ;
      RECT 0.76 0.445 0.941 0.535 ;
      RECT 2.9 0.25 2.99 0.615 ;
      RECT 1.404 0.43 1.765 0.52 ;
      RECT 1.362 0.371 1.404 0.499 ;
      RECT 1.324 0.43 1.765 0.459 ;
      RECT 0.903 0.426 1.036 0.459 ;
      RECT 0.987 0.355 0.998 0.484 ;
      RECT 0.998 0.35 1.362 0.44 ;
      RECT 1.404 0.411 1.442 0.52 ;
      RECT 0.941 0.384 0.987 0.512 ;
      RECT 2.473 0.25 2.99 0.34 ;
      RECT 2.431 0.191 2.473 0.319 ;
      RECT 2.393 0.25 2.99 0.279 ;
      RECT 2.035 0.17 2.431 0.26 ;
      RECT 2.035 0.231 2.511 0.26 ;
      RECT 0.91 0.645 1 1.01 ;
      RECT 0.225 0.72 0.315 0.86 ;
      RECT 0.225 0.72 0.542 0.81 ;
      RECT 0.225 0.72 0.617 0.754 ;
      RECT 0.58 0.645 1 0.735 ;
      RECT 0.504 0.701 1 0.735 ;
      RECT 0.542 0.663 0.58 0.791 ;
      RECT 0.58 0.215 0.67 0.735 ;
      RECT 1.855 0.25 1.945 0.6 ;
      RECT 1.48 0.25 1.945 0.34 ;
      RECT 1.438 0.191 1.48 0.319 ;
      RECT 0.58 0.215 0.915 0.305 ;
      RECT 1.4 0.25 1.945 0.279 ;
      RECT 0.825 0.17 1.438 0.26 ;
      RECT 0.58 0.231 1.518 0.26 ;
      RECT 0.045 0.945 0.185 1.035 ;
      RECT 0.045 0.28 0.135 1.035 ;
      RECT 0.045 0.515 0.49 0.605 ;
      RECT 0.4 0.465 0.49 0.605 ;
      RECT 0.045 0.28 0.185 0.37 ;
      RECT 2.55 0.93 2.92 1.02 ;
  END
END ICGNX2H7R

MACRO ICGNX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGNX3H7R 0 0 ;
  SIZE 4.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.2 1.48 ;
        RECT 3.88 1.24 4.02 1.48 ;
        RECT 3.275 1.16 3.415 1.48 ;
        RECT 2.245 1.24 2.385 1.48 ;
        RECT 1.495 1.095 1.635 1.48 ;
        RECT 0.32 1.05 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.2 0.08 ;
        RECT 3.825 -0.08 3.965 0.235 ;
        RECT 3.335 -0.08 3.425 0.36 ;
        RECT 2.55 -0.08 2.69 0.16 ;
        RECT 1.556 -0.08 1.696 0.16 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 2.45 0.51 2.79 0.6 ;
        RECT 2.625 0.455 2.79 0.6 ;
      LAYER MET2 ;
        RECT 2.65 0.23 2.75 0.76 ;
      LAYER VIA1 ;
        RECT 2.655 0.455 2.745 0.545 ;
    END
  END CKN
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.395 0.625 1.575 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END E
  PIN ECK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.855 0.325 3.945 1.069 ;
        RECT 3.54 1.065 3.901 1.114 ;
        RECT 3.799 1.046 3.945 1.069 ;
        RECT 3.837 1.018 3.855 1.146 ;
        RECT 3.585 0.325 3.945 0.415 ;
        RECT 3.54 1.065 3.837 1.155 ;
        RECT 3.585 0.255 3.675 0.415 ;
      LAYER MET2 ;
        RECT 3.85 0.23 3.95 0.76 ;
      LAYER VIA1 ;
        RECT 3.855 0.455 3.945 0.545 ;
    END
  END ECK
  OBS
    LAYER MET1 ;
      RECT 2.503 1.14 3.125 1.23 ;
      RECT 3.035 0.885 3.125 1.23 ;
      RECT 0.68 1.14 1.23 1.23 ;
      RECT 1.14 0.53 1.23 1.23 ;
      RECT 2.497 1.099 2.503 1.227 ;
      RECT 2.451 1.073 2.497 1.201 ;
      RECT 2.413 1.14 3.125 1.159 ;
      RECT 1.725 1.05 2.451 1.14 ;
      RECT 1.725 1.121 2.541 1.14 ;
      RECT 0.68 0.825 0.77 1.23 ;
      RECT 1.725 0.915 1.815 1.14 ;
      RECT 1.14 0.915 1.815 1.005 ;
      RECT 3.035 0.885 3.761 0.975 ;
      RECT 3.671 0.505 3.761 0.975 ;
      RECT 1.14 0.53 1.286 0.62 ;
      RECT 3.278 0.505 3.761 0.595 ;
      RECT 3.267 0.461 3.278 0.59 ;
      RECT 3.221 0.433 3.267 0.561 ;
      RECT 3.175 0.387 3.221 0.515 ;
      RECT 3.175 0.486 3.316 0.515 ;
      RECT 3.131 0.23 3.175 0.47 ;
      RECT 3.085 0.23 3.175 0.425 ;
      RECT 1.985 0.87 2.305 0.96 ;
      RECT 2.215 0.35 2.305 0.96 ;
      RECT 2.215 0.705 3.581 0.795 ;
      RECT 2.215 0.35 2.355 0.44 ;
      RECT 1.675 0.69 2.125 0.78 ;
      RECT 2.035 0.17 2.125 0.78 ;
      RECT 1.675 0.43 1.765 0.78 ;
      RECT 2.9 0.525 3.08 0.615 ;
      RECT 0.76 0.445 0.941 0.535 ;
      RECT 2.9 0.25 2.99 0.615 ;
      RECT 1.404 0.43 1.765 0.52 ;
      RECT 1.362 0.371 1.404 0.499 ;
      RECT 1.324 0.43 1.765 0.459 ;
      RECT 0.903 0.426 1.036 0.459 ;
      RECT 0.987 0.355 0.998 0.484 ;
      RECT 0.998 0.35 1.362 0.44 ;
      RECT 1.404 0.411 1.442 0.52 ;
      RECT 0.941 0.384 0.987 0.512 ;
      RECT 2.473 0.25 2.99 0.34 ;
      RECT 2.431 0.191 2.473 0.319 ;
      RECT 2.393 0.25 2.99 0.279 ;
      RECT 2.035 0.17 2.431 0.26 ;
      RECT 2.035 0.231 2.511 0.26 ;
      RECT 0.91 0.645 1 1.05 ;
      RECT 0.225 0.77 0.492 0.86 ;
      RECT 0.225 0.77 0.538 0.837 ;
      RECT 0.454 0.751 0.58 0.793 ;
      RECT 0.225 0.72 0.315 0.86 ;
      RECT 0.492 0.709 0.617 0.754 ;
      RECT 0.538 0.665 0.58 0.793 ;
      RECT 0.58 0.645 1 0.735 ;
      RECT 0.58 0.215 0.67 0.735 ;
      RECT 1.855 0.25 1.945 0.6 ;
      RECT 1.48 0.25 1.945 0.34 ;
      RECT 1.438 0.191 1.48 0.319 ;
      RECT 0.58 0.215 0.915 0.305 ;
      RECT 1.4 0.25 1.945 0.279 ;
      RECT 0.825 0.17 1.438 0.26 ;
      RECT 0.58 0.231 1.518 0.26 ;
      RECT 0.045 0.945 0.185 1.035 ;
      RECT 0.045 0.28 0.135 1.035 ;
      RECT 0.045 0.515 0.49 0.605 ;
      RECT 0.4 0.465 0.49 0.605 ;
      RECT 0.045 0.28 0.185 0.37 ;
      RECT 2.55 0.93 2.92 1.02 ;
  END
END ICGNX3H7R

MACRO ICGNX4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGNX4H7R 0 0 ;
  SIZE 4.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.4 1.48 ;
        RECT 3.88 1.24 4.02 1.48 ;
        RECT 3.29 1.075 3.43 1.48 ;
        RECT 2.245 1.24 2.385 1.48 ;
        RECT 1.495 1.095 1.635 1.48 ;
        RECT 0.32 1.05 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.4 0.08 ;
        RECT 3.825 -0.08 3.965 0.235 ;
        RECT 3.335 -0.08 3.425 0.36 ;
        RECT 2.55 -0.08 2.69 0.16 ;
        RECT 1.556 -0.08 1.696 0.16 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 2.45 0.51 2.79 0.6 ;
        RECT 2.625 0.455 2.79 0.6 ;
      LAYER MET2 ;
        RECT 2.65 0.23 2.75 0.76 ;
      LAYER VIA1 ;
        RECT 2.655 0.455 2.745 0.545 ;
    END
  END CKN
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.395 0.62 1.545 0.8 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END E
  PIN ECK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.855 0.952 4.3 1.042 ;
        RECT 3.855 0.325 3.945 1.042 ;
        RECT 3.855 0.325 3.941 1.071 ;
        RECT 3.54 1.065 3.901 1.114 ;
        RECT 3.799 1.046 3.941 1.071 ;
        RECT 3.837 1.018 3.855 1.146 ;
        RECT 3.56 0.325 3.945 0.415 ;
        RECT 3.54 1.065 3.837 1.155 ;
      LAYER MET2 ;
        RECT 3.85 0.23 3.95 0.76 ;
      LAYER VIA1 ;
        RECT 3.855 0.455 3.945 0.545 ;
    END
  END ECK
  OBS
    LAYER MET1 ;
      RECT 2.503 1.14 3.125 1.23 ;
      RECT 3.035 0.885 3.125 1.23 ;
      RECT 0.68 1.14 1.23 1.23 ;
      RECT 1.14 0.53 1.23 1.23 ;
      RECT 2.497 1.099 2.503 1.227 ;
      RECT 2.451 1.073 2.497 1.201 ;
      RECT 2.413 1.14 3.125 1.159 ;
      RECT 1.725 1.05 2.451 1.14 ;
      RECT 1.725 1.121 2.541 1.14 ;
      RECT 0.68 0.825 0.77 1.23 ;
      RECT 1.725 0.915 1.815 1.14 ;
      RECT 1.14 0.915 1.815 1.005 ;
      RECT 3.035 0.885 3.761 0.975 ;
      RECT 3.671 0.505 3.761 0.975 ;
      RECT 1.14 0.53 1.286 0.62 ;
      RECT 3.278 0.505 3.761 0.595 ;
      RECT 3.267 0.461 3.278 0.59 ;
      RECT 3.221 0.433 3.267 0.561 ;
      RECT 3.175 0.387 3.221 0.515 ;
      RECT 3.175 0.486 3.316 0.515 ;
      RECT 3.131 0.23 3.175 0.47 ;
      RECT 3.085 0.23 3.175 0.425 ;
      RECT 1.985 0.87 2.305 0.96 ;
      RECT 2.215 0.35 2.305 0.96 ;
      RECT 2.215 0.705 3.581 0.795 ;
      RECT 2.215 0.35 2.355 0.44 ;
      RECT 1.675 0.69 2.125 0.78 ;
      RECT 2.035 0.17 2.125 0.78 ;
      RECT 1.675 0.43 1.765 0.78 ;
      RECT 2.9 0.525 3.08 0.615 ;
      RECT 0.76 0.395 0.9 0.535 ;
      RECT 2.9 0.25 2.99 0.615 ;
      RECT 1.404 0.43 1.765 0.52 ;
      RECT 1.362 0.371 1.404 0.499 ;
      RECT 0.76 0.395 0.991 0.485 ;
      RECT 1.324 0.43 1.765 0.459 ;
      RECT 0.76 0.395 1.036 0.459 ;
      RECT 0.998 0.35 1.362 0.44 ;
      RECT 0.76 0.411 1.442 0.44 ;
      RECT 0.953 0.376 1.404 0.44 ;
      RECT 0.991 0.353 0.998 0.482 ;
      RECT 2.473 0.25 2.99 0.34 ;
      RECT 2.431 0.191 2.473 0.319 ;
      RECT 2.393 0.25 2.99 0.279 ;
      RECT 2.035 0.17 2.431 0.26 ;
      RECT 2.035 0.231 2.511 0.26 ;
      RECT 0.91 0.645 1 1.05 ;
      RECT 0.225 0.77 0.492 0.86 ;
      RECT 0.225 0.77 0.538 0.837 ;
      RECT 0.454 0.751 0.58 0.793 ;
      RECT 0.225 0.715 0.315 0.86 ;
      RECT 0.492 0.709 0.617 0.754 ;
      RECT 0.538 0.665 0.58 0.793 ;
      RECT 0.58 0.645 1 0.735 ;
      RECT 0.58 0.215 0.67 0.735 ;
      RECT 1.855 0.25 1.945 0.6 ;
      RECT 1.48 0.25 1.945 0.34 ;
      RECT 1.438 0.191 1.48 0.319 ;
      RECT 0.58 0.215 0.915 0.305 ;
      RECT 1.4 0.25 1.945 0.279 ;
      RECT 0.825 0.17 1.438 0.26 ;
      RECT 0.58 0.231 1.518 0.26 ;
      RECT 0.045 0.945 0.185 1.035 ;
      RECT 0.045 0.23 0.135 1.035 ;
      RECT 0.4 0.465 0.49 0.605 ;
      RECT 0.045 0.465 0.49 0.555 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 2.55 0.93 2.92 1.02 ;
  END
END ICGNX4H7R

MACRO ICGX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGX0P5H7R 0 0 ;
  SIZE 4.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.4 1.48 ;
        RECT 3.445 1.18 3.585 1.48 ;
        RECT 2.35 1.24 2.49 1.48 ;
        RECT 1.665 1.24 1.805 1.48 ;
        RECT 1.155 1.225 1.295 1.48 ;
        RECT 0.085 1.055 0.175 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.4 0.08 ;
        RECT 3.48 -0.08 3.62 0.16 ;
        RECT 2.672 -0.08 2.812 0.16 ;
        RECT 1.828 -0.08 1.968 0.16 ;
        RECT 1.195 -0.08 1.335 0.16 ;
        RECT 0.06 -0.08 0.2 0.325 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 2.25 0.655 2.59 0.745 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.21 0.425 0.345 0.625 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END E
  PIN ECK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 4.025 1.055 4.24 1.145 ;
        RECT 4.15 0.274 4.24 1.145 ;
      LAYER MET2 ;
        RECT 4.05 0.84 4.15 1.22 ;
      LAYER VIA1 ;
        RECT 4.055 1.055 4.145 1.145 ;
    END
  END ECK
  OBS
    LAYER MET1 ;
      RECT 2.86 1 3.791 1.09 ;
      RECT 3.2 0.25 3.97 0.34 ;
      RECT 2.634 0.25 2.85 0.34 ;
      RECT 1.79 0.25 2.006 0.34 ;
      RECT 1.035 0.25 1.373 0.34 ;
      RECT 2.928 0.21 3.29 0.3 ;
      RECT 2.124 0.17 2.516 0.26 ;
      RECT 1.491 0.17 1.672 0.26 ;
      RECT 0.805 0.17 0.917 0.26 ;
      RECT 4.016 0.25 4.06 0.881 ;
      RECT 3.97 0.25 4.016 0.926 ;
      RECT 3.967 0.822 3.97 0.951 ;
      RECT 3.921 0.847 3.967 0.975 ;
      RECT 3.875 0.893 3.921 1.021 ;
      RECT 3.829 0.939 3.875 1.067 ;
      RECT 3.791 0.981 3.829 1.09 ;
      RECT 2.89 0.21 2.928 0.319 ;
      RECT 2.888 0.211 2.89 0.339 ;
      RECT 2.85 0.231 2.888 0.34 ;
      RECT 2.596 0.231 2.634 0.34 ;
      RECT 2.554 0.191 2.596 0.319 ;
      RECT 2.516 0.17 2.554 0.279 ;
      RECT 2.086 0.17 2.124 0.279 ;
      RECT 2.044 0.191 2.086 0.319 ;
      RECT 2.006 0.231 2.044 0.34 ;
      RECT 1.752 0.231 1.79 0.34 ;
      RECT 1.71 0.191 1.752 0.319 ;
      RECT 1.672 0.17 1.71 0.279 ;
      RECT 1.453 0.17 1.491 0.279 ;
      RECT 1.411 0.191 1.453 0.319 ;
      RECT 1.373 0.231 1.411 0.34 ;
      RECT 0.997 0.231 1.035 0.34 ;
      RECT 0.955 0.191 0.997 0.319 ;
      RECT 0.917 0.17 0.955 0.279 ;
      RECT 0.445 1.14 0.91 1.23 ;
      RECT 0.82 1.045 0.91 1.23 ;
      RECT 1.457 1.06 2.745 1.15 ;
      RECT 1.442 1.06 2.745 1.143 ;
      RECT 0.445 0.485 0.535 1.23 ;
      RECT 0.82 1.045 1.48 1.135 ;
      RECT 2.655 0.878 2.745 1.15 ;
      RECT 0.82 1.052 1.495 1.135 ;
      RECT 2.655 0.878 2.766 0.929 ;
      RECT 2.655 0.878 2.804 0.899 ;
      RECT 2.701 0.833 3.779 0.88 ;
      RECT 2.745 0.8 3.836 0.846 ;
      RECT 3.779 0.746 3.79 0.875 ;
      RECT 3.79 0.43 3.88 0.801 ;
      RECT 2.766 0.79 3.88 0.801 ;
      RECT 3.741 0.771 3.779 0.88 ;
      RECT 2.97 0.43 3.88 0.52 ;
      RECT 2.97 0.39 3.11 0.52 ;
      RECT 2 0.88 2.14 0.97 ;
      RECT 2 0.475 2.09 0.97 ;
      RECT 2.877 0.61 3.7 0.7 ;
      RECT 2.872 0.569 2.877 0.698 ;
      RECT 2.826 0.544 2.872 0.672 ;
      RECT 2.78 0.498 2.826 0.626 ;
      RECT 2.78 0.591 2.915 0.626 ;
      RECT 2.742 0.475 2.78 0.584 ;
      RECT 2 0.475 2.78 0.565 ;
      RECT 2.335 0.35 2.475 0.565 ;
      RECT 1.04 0.85 1.65 0.94 ;
      RECT 1.56 0.37 1.65 0.94 ;
      RECT 1.04 0.745 1.18 0.94 ;
      RECT 1.56 0.615 1.91 0.705 ;
      RECT 1.509 0.37 1.65 0.46 ;
      RECT 0.625 0.35 0.715 1.03 ;
      RECT 1.345 0.536 1.435 0.7 ;
      RECT 1.024 0.536 1.435 0.626 ;
      RECT 1.014 0.493 1.024 0.621 ;
      RECT 0.968 0.465 1.014 0.593 ;
      RECT 0.922 0.419 0.968 0.547 ;
      RECT 0.922 0.517 1.062 0.547 ;
      RECT 0.876 0.373 0.922 0.501 ;
      RECT 0.838 0.419 0.968 0.459 ;
      RECT 0.625 0.35 0.876 0.44 ;
  END
END ICGX0P5H7R

MACRO ICGX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGX1H7R 0 0 ;
  SIZE 4.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.4 1.48 ;
        RECT 3.385 1.2 3.525 1.48 ;
        RECT 2.29 1.24 2.43 1.48 ;
        RECT 1.665 1.24 1.805 1.48 ;
        RECT 1.155 1.225 1.295 1.48 ;
        RECT 0.06 1.06 0.2 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.4 0.08 ;
        RECT 3.42 -0.08 3.56 0.16 ;
        RECT 2.612 -0.08 2.752 0.16 ;
        RECT 1.768 -0.08 1.908 0.16 ;
        RECT 1.115 -0.08 1.255 0.16 ;
        RECT 0.06 -0.08 0.2 0.325 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 2.19 0.655 2.53 0.745 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.21 0.425 0.345 0.625 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END E
  PIN ECK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 4.025 1.055 4.18 1.145 ;
        RECT 4.09 0.294 4.18 1.145 ;
      LAYER MET2 ;
        RECT 4.05 0.84 4.15 1.22 ;
      LAYER VIA1 ;
        RECT 4.055 1.055 4.145 1.145 ;
    END
  END ECK
  OBS
    LAYER MET1 ;
      RECT 2.905 1.02 3.715 1.11 ;
      RECT 3.14 0.25 3.91 0.34 ;
      RECT 2.574 0.25 2.79 0.34 ;
      RECT 1.73 0.25 1.976 0.34 ;
      RECT 1.05 0.25 1.298 0.34 ;
      RECT 2.908 0.17 3.23 0.26 ;
      RECT 2.094 0.17 2.456 0.26 ;
      RECT 1.416 0.17 1.612 0.26 ;
      RECT 0.715 0.17 0.932 0.26 ;
      RECT 3.956 0.25 4 0.885 ;
      RECT 3.91 0.25 3.956 0.93 ;
      RECT 3.891 0.834 3.91 0.963 ;
      RECT 3.845 0.867 3.891 0.995 ;
      RECT 3.799 0.913 3.845 1.041 ;
      RECT 3.753 0.959 3.799 1.087 ;
      RECT 3.715 1.001 3.753 1.11 ;
      RECT 2.87 0.17 2.908 0.279 ;
      RECT 2.828 0.191 2.87 0.319 ;
      RECT 2.79 0.231 2.828 0.34 ;
      RECT 2.536 0.231 2.574 0.34 ;
      RECT 2.494 0.191 2.536 0.319 ;
      RECT 2.456 0.17 2.494 0.279 ;
      RECT 2.056 0.17 2.094 0.279 ;
      RECT 2.014 0.191 2.056 0.319 ;
      RECT 1.976 0.231 2.014 0.34 ;
      RECT 1.692 0.231 1.73 0.34 ;
      RECT 1.65 0.191 1.692 0.319 ;
      RECT 1.612 0.17 1.65 0.279 ;
      RECT 1.378 0.17 1.416 0.279 ;
      RECT 1.336 0.191 1.378 0.319 ;
      RECT 1.298 0.231 1.336 0.34 ;
      RECT 1.012 0.231 1.05 0.34 ;
      RECT 0.97 0.191 1.012 0.319 ;
      RECT 0.932 0.17 0.97 0.279 ;
      RECT 0.445 1.14 0.92 1.23 ;
      RECT 0.83 1.045 0.92 1.23 ;
      RECT 1.457 1.06 2.686 1.15 ;
      RECT 1.442 1.06 2.686 1.143 ;
      RECT 0.445 0.485 0.535 1.23 ;
      RECT 0.83 1.045 1.48 1.135 ;
      RECT 2.596 0.848 2.686 1.15 ;
      RECT 0.83 1.052 1.495 1.135 ;
      RECT 2.596 0.848 2.715 0.895 ;
      RECT 2.596 0.848 3.719 0.88 ;
      RECT 2.642 0.807 3.73 0.875 ;
      RECT 2.677 0.79 3.776 0.846 ;
      RECT 3.719 0.746 3.73 0.875 ;
      RECT 3.73 0.43 3.82 0.801 ;
      RECT 3.681 0.771 3.82 0.801 ;
      RECT 2.91 0.43 3.82 0.52 ;
      RECT 2.91 0.39 3.05 0.52 ;
      RECT 1.96 0.88 2.1 0.97 ;
      RECT 2.01 0.475 2.1 0.97 ;
      RECT 2.717 0.61 3.64 0.7 ;
      RECT 2.712 0.569 2.717 0.698 ;
      RECT 2.666 0.544 2.712 0.672 ;
      RECT 2.62 0.498 2.666 0.626 ;
      RECT 2.62 0.591 2.755 0.626 ;
      RECT 2.582 0.475 2.62 0.584 ;
      RECT 2.01 0.475 2.62 0.565 ;
      RECT 2.275 0.35 2.415 0.565 ;
      RECT 1.01 0.85 1.585 0.94 ;
      RECT 1.495 0.37 1.585 0.94 ;
      RECT 1.01 0.72 1.15 0.94 ;
      RECT 1.495 0.615 1.92 0.705 ;
      RECT 1.495 0.37 1.59 0.705 ;
      RECT 1.449 0.37 1.59 0.46 ;
      RECT 0.625 0.37 0.715 1.03 ;
      RECT 1.043 0.54 1.405 0.63 ;
      RECT 1.003 0.482 1.043 0.61 ;
      RECT 0.957 0.439 1.003 0.567 ;
      RECT 0.957 0.521 1.081 0.567 ;
      RECT 0.911 0.393 0.957 0.521 ;
      RECT 0.873 0.439 1.003 0.479 ;
      RECT 0.625 0.37 0.911 0.46 ;
  END
END ICGX1H7R

MACRO ICGX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGX2H7R 0 0 ;
  SIZE 4.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.6 1.48 ;
        RECT 3.544 1.24 3.684 1.48 ;
        RECT 2.393 1.24 2.533 1.48 ;
        RECT 1.795 1.24 1.935 1.48 ;
        RECT 1.255 1.225 1.395 1.48 ;
        RECT 0.06 1.06 0.2 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.6 0.08 ;
        RECT 3.534 -0.08 3.674 0.16 ;
        RECT 2.712 -0.08 2.852 0.16 ;
        RECT 1.873 -0.08 2.013 0.16 ;
        RECT 1.245 -0.08 1.385 0.16 ;
        RECT 0.06 -0.08 0.2 0.325 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 2.332 0.745 2.672 0.945 ;
      LAYER MET2 ;
        RECT 2.45 0.625 2.55 1.16 ;
      LAYER VIA1 ;
        RECT 2.455 0.855 2.545 0.945 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.21 0.425 0.345 0.625 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END E
  PIN ECK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 4.204 1.025 4.345 1.175 ;
        RECT 4.204 0.229 4.294 1.175 ;
      LAYER MET2 ;
        RECT 4.25 0.84 4.35 1.22 ;
      LAYER VIA1 ;
        RECT 4.255 1.055 4.345 1.145 ;
    END
  END ECK
  OBS
    LAYER MET1 ;
      RECT 2.966 1.06 4.114 1.15 ;
      RECT 4.024 0.25 4.114 1.15 ;
      RECT 3.239 0.25 4.114 0.34 ;
      RECT 2.636 0.25 2.928 0.34 ;
      RECT 1.797 0.25 2.104 0.34 ;
      RECT 1.167 0.25 1.461 0.34 ;
      RECT 2.594 0.25 2.97 0.319 ;
      RECT 1.755 0.25 2.146 0.319 ;
      RECT 1.125 0.25 1.503 0.319 ;
      RECT 2.556 0.25 3.008 0.279 ;
      RECT 1.717 0.25 2.184 0.279 ;
      RECT 1.087 0.25 1.541 0.279 ;
      RECT 2.97 0.17 3.329 0.26 ;
      RECT 2.89 0.231 3.329 0.26 ;
      RECT 2.928 0.191 2.97 0.319 ;
      RECT 2.066 0.231 2.674 0.26 ;
      RECT 1.423 0.231 1.835 0.26 ;
      RECT 0.805 0.231 1.205 0.26 ;
      RECT 2.104 0.191 2.636 0.26 ;
      RECT 1.461 0.191 1.797 0.26 ;
      RECT 0.805 0.191 1.167 0.26 ;
      RECT 2.146 0.17 2.594 0.26 ;
      RECT 1.503 0.17 1.755 0.26 ;
      RECT 0.805 0.17 1.125 0.26 ;
      RECT 0.445 1.14 0.985 1.23 ;
      RECT 0.895 1.045 0.985 1.23 ;
      RECT 1.457 1.06 2.851 1.15 ;
      RECT 1.442 1.06 2.851 1.143 ;
      RECT 0.445 0.485 0.535 1.23 ;
      RECT 0.895 1.045 1.48 1.135 ;
      RECT 2.761 0.979 2.851 1.15 ;
      RECT 0.895 1.052 1.495 1.135 ;
      RECT 2.807 0.934 2.897 1.017 ;
      RECT 2.851 0.889 2.943 0.971 ;
      RECT 2.897 0.843 3.011 0.899 ;
      RECT 2.943 0.805 2.973 0.933 ;
      RECT 3.844 0.43 3.934 0.88 ;
      RECT 2.973 0.79 3.934 0.88 ;
      RECT 3.009 0.43 3.934 0.52 ;
      RECT 3.009 0.39 3.149 0.52 ;
      RECT 2.09 0.565 2.23 0.97 ;
      RECT 2.802 0.61 3.754 0.7 ;
      RECT 2.795 0.568 2.802 0.697 ;
      RECT 2.757 0.61 3.754 0.674 ;
      RECT 2.09 0.565 2.795 0.655 ;
      RECT 2.09 0.591 2.84 0.655 ;
      RECT 2.37 0.35 2.518 0.655 ;
      RECT 1.04 0.85 1.699 0.94 ;
      RECT 1.559 0.37 1.699 0.94 ;
      RECT 1.04 0.745 1.18 0.94 ;
      RECT 1.559 0.615 1.967 0.705 ;
      RECT 0.625 0.35 0.715 1.03 ;
      RECT 1.36 0.536 1.45 0.7 ;
      RECT 1.194 0.536 1.45 0.626 ;
      RECT 1.184 0.493 1.194 0.621 ;
      RECT 1.138 0.465 1.184 0.593 ;
      RECT 1.092 0.419 1.138 0.547 ;
      RECT 1.092 0.517 1.232 0.547 ;
      RECT 1.046 0.373 1.092 0.501 ;
      RECT 1.008 0.419 1.138 0.459 ;
      RECT 0.625 0.35 1.046 0.44 ;
  END
END ICGX2H7R

MACRO ICGX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGX3H7R 0 0 ;
  SIZE 4.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.8 1.48 ;
        RECT 4.454 0.99 4.544 1.48 ;
        RECT 3.544 1.24 3.684 1.48 ;
        RECT 2.412 1.24 2.552 1.48 ;
        RECT 1.795 1.24 1.935 1.48 ;
        RECT 1.255 1.225 1.395 1.48 ;
        RECT 0.06 1.06 0.2 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.8 0.08 ;
        RECT 4.454 -0.08 4.544 0.355 ;
        RECT 3.55 -0.08 3.69 0.16 ;
        RECT 2.745 -0.08 2.885 0.16 ;
        RECT 1.873 -0.08 2.013 0.16 ;
        RECT 1.245 -0.08 1.385 0.16 ;
        RECT 0.06 -0.08 0.2 0.325 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 2.332 0.745 2.672 0.945 ;
      LAYER MET2 ;
        RECT 2.45 0.625 2.55 1.16 ;
      LAYER VIA1 ;
        RECT 2.455 0.855 2.545 0.945 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.21 0.425 0.345 0.625 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END E
  PIN ECK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 4.204 0.825 4.345 1.035 ;
        RECT 4.204 0.229 4.294 1.035 ;
      LAYER MET2 ;
        RECT 4.25 0.625 4.35 1.16 ;
      LAYER VIA1 ;
        RECT 4.255 0.855 4.345 0.945 ;
    END
  END ECK
  OBS
    LAYER MET1 ;
      RECT 2.966 1.06 4.114 1.15 ;
      RECT 4.024 0.25 4.114 1.15 ;
      RECT 3.27 0.25 4.114 0.34 ;
      RECT 2.669 0.25 2.961 0.34 ;
      RECT 1.797 0.25 2.104 0.34 ;
      RECT 1.167 0.25 1.461 0.34 ;
      RECT 2.627 0.25 3.003 0.319 ;
      RECT 1.755 0.25 2.146 0.319 ;
      RECT 1.125 0.25 1.503 0.319 ;
      RECT 2.589 0.25 3.041 0.279 ;
      RECT 1.717 0.25 2.184 0.279 ;
      RECT 1.087 0.25 1.541 0.279 ;
      RECT 3.003 0.17 3.36 0.26 ;
      RECT 2.923 0.231 3.36 0.26 ;
      RECT 2.961 0.191 3.003 0.319 ;
      RECT 2.066 0.231 2.707 0.26 ;
      RECT 1.423 0.231 1.835 0.26 ;
      RECT 0.805 0.231 1.205 0.26 ;
      RECT 2.104 0.191 2.669 0.26 ;
      RECT 1.461 0.191 1.797 0.26 ;
      RECT 0.805 0.191 1.167 0.26 ;
      RECT 2.146 0.17 2.627 0.26 ;
      RECT 1.503 0.17 1.755 0.26 ;
      RECT 0.805 0.17 1.125 0.26 ;
      RECT 0.445 1.14 0.985 1.23 ;
      RECT 0.895 1.045 0.985 1.23 ;
      RECT 1.457 1.06 2.851 1.15 ;
      RECT 1.442 1.06 2.851 1.143 ;
      RECT 0.445 0.485 0.535 1.23 ;
      RECT 0.895 1.045 1.48 1.135 ;
      RECT 2.761 0.979 2.851 1.15 ;
      RECT 0.895 1.052 1.495 1.135 ;
      RECT 2.807 0.934 2.897 1.017 ;
      RECT 2.851 0.889 2.943 0.971 ;
      RECT 2.897 0.843 3.011 0.899 ;
      RECT 2.943 0.805 2.973 0.933 ;
      RECT 3.844 0.43 3.934 0.88 ;
      RECT 2.973 0.79 3.934 0.88 ;
      RECT 3.04 0.43 3.934 0.52 ;
      RECT 3.04 0.39 3.18 0.52 ;
      RECT 2.09 0.565 2.23 0.97 ;
      RECT 2.802 0.61 3.754 0.7 ;
      RECT 2.795 0.568 2.802 0.697 ;
      RECT 2.757 0.61 3.754 0.674 ;
      RECT 2.09 0.565 2.795 0.655 ;
      RECT 2.09 0.591 2.84 0.655 ;
      RECT 2.413 0.36 2.561 0.655 ;
      RECT 1.04 0.85 1.699 0.94 ;
      RECT 1.559 0.37 1.699 0.94 ;
      RECT 1.04 0.745 1.18 0.94 ;
      RECT 1.559 0.615 1.967 0.705 ;
      RECT 0.625 0.35 0.715 1.03 ;
      RECT 1.36 0.536 1.45 0.7 ;
      RECT 1.194 0.536 1.45 0.626 ;
      RECT 1.184 0.493 1.194 0.621 ;
      RECT 1.138 0.465 1.184 0.593 ;
      RECT 1.092 0.419 1.138 0.547 ;
      RECT 1.092 0.517 1.232 0.547 ;
      RECT 1.046 0.373 1.092 0.501 ;
      RECT 1.008 0.419 1.138 0.459 ;
      RECT 0.625 0.35 1.046 0.44 ;
  END
END ICGX3H7R

MACRO ICGX4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICGX4H7R 0 0 ;
  SIZE 4.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.8 1.48 ;
        RECT 4.454 0.99 4.544 1.48 ;
        RECT 3.544 1.24 3.684 1.48 ;
        RECT 2.412 1.24 2.552 1.48 ;
        RECT 1.795 1.24 1.935 1.48 ;
        RECT 1.255 1.225 1.395 1.48 ;
        RECT 0.06 1.06 0.2 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.8 0.08 ;
        RECT 4.44 -0.08 4.53 0.355 ;
        RECT 3.55 -0.08 3.69 0.16 ;
        RECT 2.745 -0.08 2.885 0.16 ;
        RECT 1.873 -0.08 2.013 0.16 ;
        RECT 1.245 -0.08 1.385 0.16 ;
        RECT 0.06 -0.08 0.2 0.325 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 2.332 0.745 2.672 0.945 ;
      LAYER MET2 ;
        RECT 2.45 0.625 2.55 1.16 ;
      LAYER VIA1 ;
        RECT 2.455 0.855 2.545 0.945 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.21 0.425 0.345 0.625 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END E
  PIN ECK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 4.19 1.025 4.345 1.175 ;
        RECT 4.19 0.349 4.28 1.175 ;
      LAYER MET2 ;
        RECT 4.25 0.84 4.35 1.22 ;
      LAYER VIA1 ;
        RECT 4.255 1.055 4.345 1.145 ;
    END
  END ECK
  OBS
    LAYER MET1 ;
      RECT 2.966 1.06 4.1 1.15 ;
      RECT 4.01 0.25 4.1 1.15 ;
      RECT 3.27 0.25 4.1 0.34 ;
      RECT 2.669 0.25 2.961 0.34 ;
      RECT 1.797 0.25 2.104 0.34 ;
      RECT 1.167 0.25 1.461 0.34 ;
      RECT 2.627 0.25 3.003 0.319 ;
      RECT 1.755 0.25 2.146 0.319 ;
      RECT 1.125 0.25 1.503 0.319 ;
      RECT 2.589 0.25 3.041 0.279 ;
      RECT 1.717 0.25 2.184 0.279 ;
      RECT 1.087 0.25 1.541 0.279 ;
      RECT 3.003 0.17 3.36 0.26 ;
      RECT 2.923 0.231 3.36 0.26 ;
      RECT 2.961 0.191 3.003 0.319 ;
      RECT 2.066 0.231 2.707 0.26 ;
      RECT 1.423 0.231 1.835 0.26 ;
      RECT 0.805 0.231 1.205 0.26 ;
      RECT 2.104 0.191 2.669 0.26 ;
      RECT 1.461 0.191 1.797 0.26 ;
      RECT 0.805 0.191 1.167 0.26 ;
      RECT 2.146 0.17 2.627 0.26 ;
      RECT 1.503 0.17 1.755 0.26 ;
      RECT 0.805 0.17 1.125 0.26 ;
      RECT 0.445 1.14 0.985 1.23 ;
      RECT 0.895 1.045 0.985 1.23 ;
      RECT 1.457 1.06 2.851 1.15 ;
      RECT 1.442 1.06 2.851 1.143 ;
      RECT 0.445 0.485 0.535 1.23 ;
      RECT 0.895 1.045 1.48 1.135 ;
      RECT 2.761 0.979 2.851 1.15 ;
      RECT 0.895 1.052 1.495 1.135 ;
      RECT 2.807 0.934 2.897 1.017 ;
      RECT 2.851 0.889 2.943 0.971 ;
      RECT 2.897 0.843 3.011 0.899 ;
      RECT 2.943 0.805 2.973 0.933 ;
      RECT 3.83 0.43 3.92 0.88 ;
      RECT 2.973 0.79 3.92 0.88 ;
      RECT 3.04 0.43 3.92 0.52 ;
      RECT 3.04 0.39 3.18 0.52 ;
      RECT 2.09 0.565 2.23 0.97 ;
      RECT 2.802 0.61 3.74 0.7 ;
      RECT 2.795 0.568 2.802 0.697 ;
      RECT 2.757 0.61 3.74 0.674 ;
      RECT 2.09 0.565 2.795 0.655 ;
      RECT 2.09 0.591 2.84 0.655 ;
      RECT 2.413 0.36 2.561 0.655 ;
      RECT 1.04 0.85 1.699 0.94 ;
      RECT 1.559 0.37 1.699 0.94 ;
      RECT 1.04 0.745 1.18 0.94 ;
      RECT 1.559 0.615 1.967 0.705 ;
      RECT 0.625 0.35 0.715 1.03 ;
      RECT 1.36 0.536 1.45 0.7 ;
      RECT 1.194 0.536 1.45 0.626 ;
      RECT 1.184 0.493 1.194 0.621 ;
      RECT 1.138 0.465 1.184 0.593 ;
      RECT 1.092 0.419 1.138 0.547 ;
      RECT 1.092 0.517 1.232 0.547 ;
      RECT 1.046 0.373 1.092 0.501 ;
      RECT 1.008 0.419 1.138 0.459 ;
      RECT 0.625 0.35 1.046 0.44 ;
  END
END ICGX4H7R

MACRO INVX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX0P5H7R 0 0 ;
  SIZE 0.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.6 1.48 ;
        RECT 0.07 1 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.6 0.08 ;
        RECT 0.07 -0.08 0.16 0.45 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.165 0.625 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.305 1.015 0.545 1.105 ;
        RECT 0.455 0.335 0.545 1.105 ;
        RECT 0.315 0.335 0.545 0.425 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END Y
END INVX0P5H7R

MACRO INVX0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX0P7H7R 0 0 ;
  SIZE 0.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.6 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.6 0.08 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.05 0.625 0.23 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.32 0.225 0.545 0.375 ;
        RECT 0.32 0.225 0.41 1.123 ;
      LAYER MET2 ;
        RECT 0.45 0.18 0.55 0.56 ;
      LAYER VIA1 ;
        RECT 0.455 0.255 0.545 0.345 ;
    END
  END Y
END INVX0P7H7R

MACRO INVX10H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX10H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.07 1.07 1.16 1.48 ;
        RECT 0.57 1.07 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.57 -0.08 1.66 0.345 ;
        RECT 1.07 -0.08 1.16 0.33 ;
        RECT 0.57 -0.08 0.66 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.655 1.19 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.295 0.885 1.41 0.975 ;
        RECT 1.32 0.22 1.41 0.975 ;
        RECT 0.32 0.455 1.41 0.545 ;
        RECT 0.82 0.37 0.91 0.545 ;
        RECT 0.32 0.22 0.41 0.545 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END Y
END INVX10H7R

MACRO INVX12H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX12H7R 0 0 ;
  SIZE 3.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.4 1.48 ;
        RECT 3.235 1.05 3.325 1.48 ;
        RECT 2.705 1.05 2.795 1.48 ;
        RECT 2.175 1.05 2.265 1.48 ;
        RECT 1.645 1.05 1.735 1.48 ;
        RECT 1.115 1.05 1.205 1.48 ;
        RECT 0.585 1.05 0.675 1.48 ;
        RECT 0.07 0.905 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.4 0.08 ;
        RECT 3.235 -0.08 3.325 0.235 ;
        RECT 2.705 -0.08 2.795 0.235 ;
        RECT 2.175 -0.08 2.265 0.235 ;
        RECT 1.645 -0.08 1.735 0.235 ;
        RECT 1.115 -0.08 1.205 0.235 ;
        RECT 0.585 -0.08 0.675 0.235 ;
        RECT 0.07 -0.08 0.16 0.45 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.615 3.135 0.705 ;
        RECT 0.055 0.615 0.145 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.32 0.805 3.345 0.895 ;
        RECT 3.255 0.335 3.345 0.895 ;
        RECT 0.295 0.335 3.345 0.425 ;
        RECT 2.97 0.805 3.06 1.045 ;
        RECT 2.44 0.805 2.53 1.045 ;
        RECT 1.91 0.805 2 1.045 ;
        RECT 1.38 0.805 1.47 1.045 ;
        RECT 0.85 0.805 0.94 1.045 ;
        RECT 0.32 0.805 0.41 1.045 ;
      LAYER MET2 ;
        RECT 3.25 0.23 3.35 0.76 ;
      LAYER VIA1 ;
        RECT 3.255 0.455 3.345 0.545 ;
    END
  END Y
END INVX12H7R

MACRO INVX16H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX16H7R 0 0 ;
  SIZE 3.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.6 1.48 ;
        RECT 2.97 1 3.06 1.48 ;
        RECT 2.77 1 3.06 1.14 ;
        RECT 2.07 1 2.16 1.48 ;
        RECT 1.87 1 2.16 1.155 ;
        RECT 1.17 1 1.26 1.48 ;
        RECT 0.97 1 1.26 1.14 ;
        RECT 0.27 0.8 0.36 1.48 ;
        RECT 0.07 0.8 0.36 1.14 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.6 0.08 ;
        RECT 3.045 -0.08 3.185 0.305 ;
        RECT 2.545 -0.08 2.685 0.305 ;
        RECT 2.045 -0.08 2.185 0.305 ;
        RECT 1.545 -0.08 1.685 0.305 ;
        RECT 1.045 -0.08 1.185 0.305 ;
        RECT 0.545 -0.08 0.685 0.305 ;
        RECT 0.045 -0.08 0.185 0.32 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.575 3.165 0.665 ;
        RECT 0.055 0.425 0.145 0.665 ;
      LAYER MET2 ;
        RECT 0.05 0.23 0.15 0.76 ;
      LAYER VIA1 ;
        RECT 0.055 0.455 0.145 0.545 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.22 1 3.51 1.145 ;
        RECT 3.42 0.26 3.51 1.145 ;
        RECT 0.72 0.755 3.51 0.845 ;
        RECT 0.32 0.395 3.51 0.485 ;
        RECT 2.82 0.265 2.91 0.485 ;
        RECT 2.32 1 2.61 1.14 ;
        RECT 2.52 0.755 2.61 1.14 ;
        RECT 2.32 0.265 2.41 0.485 ;
        RECT 1.82 0.265 1.91 0.485 ;
        RECT 1.42 1 1.71 1.14 ;
        RECT 1.62 0.755 1.71 1.14 ;
        RECT 1.32 0.265 1.41 0.485 ;
        RECT 0.82 0.265 0.91 0.485 ;
        RECT 0.52 1 0.81 1.14 ;
        RECT 0.72 0.755 0.81 1.14 ;
        RECT 0.32 0.265 0.41 0.485 ;
      LAYER MET2 ;
        RECT 3.25 0.84 3.35 1.22 ;
      LAYER VIA1 ;
        RECT 3.255 1.055 3.345 1.145 ;
    END
  END Y
END INVX16H7R

MACRO INVX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX1H7R 0 0 ;
  SIZE 0.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.6 1.48 ;
        RECT 0.07 1.02 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.6 0.08 ;
        RECT 0.07 -0.08 0.16 0.39 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.305 0.925 0.545 1.015 ;
        RECT 0.455 0.335 0.545 1.015 ;
        RECT 0.315 0.335 0.545 0.425 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END Y
END INVX1H7R

MACRO INVX1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX1P4H7R 0 0 ;
  SIZE 0.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.6 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.6 0.08 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.05 0.625 0.23 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.32 0.225 0.41 1.031 ;
        RECT 0.255 0.225 0.41 0.375 ;
      LAYER MET2 ;
        RECT 0.25 0.18 0.35 0.56 ;
      LAYER VIA1 ;
        RECT 0.255 0.255 0.345 0.345 ;
    END
  END Y
END INVX1P4H7R

MACRO INVX20H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX20H7R 0 0 ;
  SIZE 3 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3 1.48 ;
        RECT 2.57 1.055 2.66 1.48 ;
        RECT 2.07 1.07 2.16 1.48 ;
        RECT 1.57 1.07 1.66 1.48 ;
        RECT 1.07 1.07 1.16 1.48 ;
        RECT 0.57 1.07 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3 0.08 ;
        RECT 2.57 -0.08 2.66 0.33 ;
        RECT 2.045 -0.08 2.185 0.305 ;
        RECT 1.545 -0.08 1.685 0.305 ;
        RECT 1.045 -0.08 1.185 0.305 ;
        RECT 0.545 -0.08 0.685 0.305 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.655 2.19 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.345 0.455 2.91 0.545 ;
        RECT 2.82 0.205 2.91 0.545 ;
        RECT 0.295 0.885 2.435 0.975 ;
        RECT 2.345 0.395 2.435 0.975 ;
        RECT 0.32 0.395 2.435 0.485 ;
        RECT 0.32 0.22 0.41 0.485 ;
      LAYER MET2 ;
        RECT 2.65 0.23 2.75 0.76 ;
      LAYER VIA1 ;
        RECT 2.655 0.455 2.745 0.545 ;
    END
  END Y
END INVX20H7R

MACRO INVX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX2H7R 0 0 ;
  SIZE 0.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.8 1.48 ;
        RECT 0.63 1.055 0.72 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.8 0.08 ;
        RECT 0.63 -0.08 0.72 0.38 ;
        RECT 0.07 -0.08 0.16 0.38 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.22 0.655 0.565 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.32 0.875 0.745 0.965 ;
        RECT 0.655 0.47 0.745 0.965 ;
        RECT 0.35 0.47 0.745 0.56 ;
        RECT 0.35 0.24 0.44 0.56 ;
        RECT 0.32 0.875 0.41 1.2 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END Y
END INVX2H7R

MACRO INVX2P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX2P5H7R 0 0 ;
  SIZE 0.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.8 1.48 ;
        RECT 0.57 1.055 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.8 0.08 ;
        RECT 0.57 -0.08 0.66 0.345 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.05 0.625 0.23 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.32 0.225 0.41 1.095 ;
        RECT 0.255 0.225 0.41 0.375 ;
      LAYER MET2 ;
        RECT 0.25 0.18 0.35 0.56 ;
      LAYER VIA1 ;
        RECT 0.255 0.255 0.345 0.345 ;
    END
  END Y
END INVX2P5H7R

MACRO INVX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX3H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.58 1.03 0.67 1.48 ;
        RECT 0.07 1.03 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.555 -0.08 0.695 0.365 ;
        RECT 0.07 -0.08 0.16 0.39 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.655 0.765 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.84 0.85 0.945 1.17 ;
        RECT 0.855 0.455 0.945 1.17 ;
        RECT 0.32 0.455 0.945 0.545 ;
        RECT 0.32 0.85 0.945 0.94 ;
        RECT 0.32 0.85 0.41 1.17 ;
        RECT 0.32 0.25 0.41 0.545 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
END INVX3H7R

MACRO INVX3P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX3P5H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.57 1.055 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.57 -0.08 0.66 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.05 0.625 0.23 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.32 0.455 0.91 0.545 ;
        RECT 0.82 0.23 0.91 0.545 ;
        RECT 0.32 0.245 0.41 1 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END Y
END INVX3P5H7R

MACRO INVX4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX4H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.24 1.035 1.33 1.48 ;
        RECT 0.6 1.035 0.69 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.24 -0.08 1.33 0.45 ;
        RECT 0.585 -0.08 0.675 0.245 ;
        RECT 0.07 -0.08 0.16 0.45 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.655 0.965 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.32 0.855 1.145 0.945 ;
        RECT 1.055 0.335 1.145 0.945 ;
        RECT 0.295 0.335 1.145 0.425 ;
        RECT 0.85 0.855 0.94 1.175 ;
        RECT 0.32 0.855 0.41 1.175 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END Y
END INVX4H7R

MACRO INVX5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX5H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.57 1.07 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.57 -0.08 0.66 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.115 0.655 0.655 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.82 0.305 0.91 0.995 ;
        RECT 0.32 0.855 0.91 0.945 ;
        RECT 0.32 0.42 0.91 0.51 ;
        RECT 0.32 0.855 0.41 1.03 ;
        RECT 0.32 0.32 0.41 0.51 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END Y
END INVX5H7R

MACRO INVX6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX6H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.67 1.12 1.76 1.48 ;
        RECT 1.115 1.12 1.205 1.48 ;
        RECT 0.585 1.12 0.675 1.48 ;
        RECT 0.07 0.98 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.685 -0.08 1.775 0.255 ;
        RECT 1.115 -0.08 1.205 0.255 ;
        RECT 0.585 -0.08 0.675 0.255 ;
        RECT 0.07 -0.08 0.16 0.45 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.655 1.575 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.32 0.92 1.76 1.01 ;
        RECT 1.67 0.35 1.76 1.01 ;
        RECT 0.295 0.35 1.76 0.44 ;
        RECT 1.39 0.92 1.48 1.08 ;
        RECT 0.85 0.92 0.945 1.175 ;
        RECT 0.32 0.92 0.41 1.08 ;
      LAYER MET2 ;
        RECT 0.85 0.84 0.95 1.22 ;
      LAYER VIA1 ;
        RECT 0.855 1.055 0.945 1.145 ;
    END
  END Y
END INVX6H7R

MACRO INVX7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX7H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.045 1.08 1.185 1.48 ;
        RECT 0.57 1.07 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.07 -0.08 1.16 0.33 ;
        RECT 0.57 -0.08 0.66 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.29 0.655 1.23 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.295 0.885 1.41 0.975 ;
        RECT 1.32 0.205 1.41 0.975 ;
        RECT 0.32 0.455 1.41 0.545 ;
        RECT 0.82 0.37 0.91 0.545 ;
        RECT 0.32 0.22 0.41 0.545 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END Y
END INVX7H7R

MACRO INVX8H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX8H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 2.28 1.11 2.37 1.48 ;
        RECT 1.735 1.11 1.825 1.48 ;
        RECT 1.13 1.11 1.22 1.48 ;
        RECT 0.6 1.11 0.69 1.48 ;
        RECT 0.07 0.93 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 2.28 -0.08 2.37 0.245 ;
        RECT 1.735 -0.08 1.825 0.245 ;
        RECT 1.13 -0.08 1.22 0.245 ;
        RECT 0.6 -0.08 0.69 0.245 ;
        RECT 0.07 -0.08 0.16 0.45 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.655 2.165 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.295 0.92 2.345 1.01 ;
        RECT 2.255 0.335 2.345 1.01 ;
        RECT 0.295 0.335 2.345 0.425 ;
      LAYER MET2 ;
        RECT 2.25 0.23 2.35 0.76 ;
      LAYER VIA1 ;
        RECT 2.255 0.455 2.345 0.545 ;
    END
  END Y
END INVX8H7R

MACRO LATHRX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATHRX0P5H7R 0 0 ;
  SIZE 4.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.2 1.48 ;
        RECT 3.61 1.18 3.75 1.48 ;
        RECT 3.05 1.18 3.19 1.48 ;
        RECT 2.615 1.055 2.705 1.48 ;
        RECT 1.82 1.24 1.96 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.2 0.08 ;
        RECT 3.73 -0.08 3.82 0.345 ;
        RECT 3.25 -0.08 3.34 0.33 ;
        RECT 2.02 -0.08 2.16 0.16 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.655 0.562 1.745 0.777 ;
        RECT 1.57 0.562 1.745 0.652 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.455 0.375 0.635 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END G
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.455 0.28 3.615 0.37 ;
        RECT 3.315 0.82 3.545 0.91 ;
        RECT 3.455 0.28 3.545 0.91 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.825 0.855 4.07 0.945 ;
        RECT 3.98 0.255 4.07 0.945 ;
      LAYER MET2 ;
        RECT 3.85 0.63 3.95 1.16 ;
      LAYER VIA1 ;
        RECT 3.855 0.855 3.945 0.945 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.96 0.455 2.175 0.545 ;
        RECT 1.96 0.455 2.05 0.63 ;
      LAYER MET2 ;
        RECT 2.05 0.23 2.15 0.76 ;
      LAYER VIA1 ;
        RECT 2.055 0.455 2.145 0.545 ;
    END
  END RN
  OBS
    LAYER MET1 ;
      RECT 3.055 1 3.725 1.09 ;
      RECT 3.635 0.668 3.725 1.09 ;
      RECT 3.055 0.255 3.145 1.09 ;
      RECT 2.44 0.82 3.145 0.91 ;
      RECT 3.635 0.668 3.89 0.76 ;
      RECT 3.8 0.62 3.89 0.76 ;
      RECT 3 0.255 3.145 0.395 ;
      RECT 1.089 0.96 1.623 1.05 ;
      RECT 1.089 0.96 1.709 0.987 ;
      RECT 1.089 0.96 1.713 0.962 ;
      RECT 2.185 0.64 2.275 0.96 ;
      RECT 1.663 0.87 2.275 0.96 ;
      RECT 1.573 0.937 2.275 0.96 ;
      RECT 1.623 0.89 1.663 1.03 ;
      RECT 1.089 0.35 1.179 1.05 ;
      RECT 1.619 0.912 2.275 0.96 ;
      RECT 2.185 0.64 2.965 0.73 ;
      RECT 2.82 0.57 2.965 0.73 ;
      RECT 2.82 0.25 2.91 0.73 ;
      RECT 0.965 0.35 1.179 0.44 ;
      RECT 2.72 0.25 2.91 0.34 ;
      RECT 0.045 0.725 0.16 1.065 ;
      RECT 0.045 0.725 0.569 0.815 ;
      RECT 0.479 0.675 0.569 0.815 ;
      RECT 0.045 0.275 0.135 1.065 ;
      RECT 2.507 0.46 2.73 0.55 ;
      RECT 2.507 0.25 2.597 0.55 ;
      RECT 0.045 0.275 0.517 0.365 ;
      RECT 1.748 0.25 2.597 0.34 ;
      RECT 1.707 0.19 1.748 0.32 ;
      RECT 1.668 0.25 2.597 0.28 ;
      RECT 0.479 0.256 0.622 0.279 ;
      RECT 0.563 0.18 0.584 0.309 ;
      RECT 0.584 0.17 1.707 0.26 ;
      RECT 0.517 0.214 0.563 0.342 ;
      RECT 0.517 0.23 1.787 0.26 ;
      RECT 0.839 1.14 1.699 1.23 ;
      RECT 2.365 1.055 2.455 1.195 ;
      RECT 0.839 1.14 1.746 1.184 ;
      RECT 0.839 1.14 1.784 1.164 ;
      RECT 1.745 1.055 2.455 1.145 ;
      RECT 1.661 1.121 2.455 1.145 ;
      RECT 1.699 1.079 1.745 1.207 ;
      RECT 0.839 0.847 0.929 1.23 ;
      RECT 1.375 0.78 1.534 0.87 ;
      RECT 1.375 0.35 1.465 0.87 ;
      RECT 1.375 0.35 1.515 0.44 ;
      RECT 0.56 0.95 0.749 1.04 ;
      RECT 0.659 0.645 0.749 1.04 ;
      RECT 0.659 0.645 0.845 0.735 ;
      RECT 0.755 0.35 0.845 0.735 ;
      RECT 0.66 0.35 0.845 0.44 ;
  END
END LATHRX0P5H7R

MACRO LATHRX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATHRX1H7R 0 0 ;
  SIZE 4.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.2 1.48 ;
        RECT 3.62 1.18 3.76 1.48 ;
        RECT 3.05 1.18 3.19 1.48 ;
        RECT 2.615 1.055 2.705 1.48 ;
        RECT 1.82 1.24 1.96 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.2 0.08 ;
        RECT 3.75 -0.08 3.84 0.345 ;
        RECT 3.25 -0.08 3.34 0.33 ;
        RECT 2.02 -0.08 2.16 0.16 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.655 0.562 1.745 0.777 ;
        RECT 1.57 0.562 1.745 0.652 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.455 0.375 0.635 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END G
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.455 0.32 3.615 0.41 ;
        RECT 3.315 0.82 3.545 0.91 ;
        RECT 3.455 0.32 3.545 0.91 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.825 0.855 4.11 0.945 ;
        RECT 4.02 0.295 4.11 0.945 ;
      LAYER MET2 ;
        RECT 3.85 0.63 3.95 1.16 ;
      LAYER VIA1 ;
        RECT 3.855 0.855 3.945 0.945 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.96 0.455 2.175 0.545 ;
        RECT 1.96 0.455 2.05 0.63 ;
      LAYER MET2 ;
        RECT 2.05 0.23 2.15 0.76 ;
      LAYER VIA1 ;
        RECT 2.055 0.455 2.145 0.545 ;
    END
  END RN
  OBS
    LAYER MET1 ;
      RECT 3.055 1 3.725 1.09 ;
      RECT 3.635 0.668 3.725 1.09 ;
      RECT 3.055 0.255 3.145 1.09 ;
      RECT 2.44 0.82 3.145 0.91 ;
      RECT 3.635 0.668 3.93 0.76 ;
      RECT 3.84 0.62 3.93 0.76 ;
      RECT 3 0.255 3.145 0.395 ;
      RECT 1.089 0.96 1.623 1.05 ;
      RECT 1.089 0.96 1.709 0.987 ;
      RECT 1.089 0.96 1.713 0.962 ;
      RECT 2.185 0.64 2.275 0.96 ;
      RECT 1.663 0.87 2.275 0.96 ;
      RECT 1.573 0.937 2.275 0.96 ;
      RECT 1.623 0.89 1.663 1.03 ;
      RECT 1.089 0.35 1.179 1.05 ;
      RECT 1.619 0.912 2.275 0.96 ;
      RECT 2.185 0.64 2.965 0.73 ;
      RECT 2.82 0.57 2.965 0.73 ;
      RECT 2.82 0.25 2.91 0.73 ;
      RECT 0.965 0.35 1.179 0.44 ;
      RECT 2.72 0.25 2.91 0.34 ;
      RECT 0.045 0.725 0.16 1.065 ;
      RECT 0.045 0.725 0.569 0.815 ;
      RECT 0.479 0.675 0.569 0.815 ;
      RECT 0.045 0.275 0.135 1.065 ;
      RECT 2.507 0.46 2.73 0.55 ;
      RECT 2.507 0.25 2.597 0.55 ;
      RECT 0.045 0.275 0.517 0.365 ;
      RECT 1.748 0.25 2.597 0.34 ;
      RECT 1.707 0.19 1.748 0.32 ;
      RECT 1.668 0.25 2.597 0.28 ;
      RECT 0.479 0.256 0.622 0.279 ;
      RECT 0.563 0.18 0.584 0.309 ;
      RECT 0.584 0.17 1.707 0.26 ;
      RECT 0.517 0.214 0.563 0.342 ;
      RECT 0.517 0.23 1.787 0.26 ;
      RECT 0.839 1.14 1.699 1.23 ;
      RECT 2.365 1.055 2.455 1.195 ;
      RECT 0.839 1.14 1.746 1.184 ;
      RECT 0.839 1.14 1.784 1.164 ;
      RECT 1.745 1.055 2.455 1.145 ;
      RECT 1.661 1.121 2.455 1.145 ;
      RECT 1.699 1.079 1.745 1.207 ;
      RECT 0.839 0.847 0.929 1.23 ;
      RECT 1.375 0.78 1.534 0.87 ;
      RECT 1.375 0.35 1.465 0.87 ;
      RECT 1.375 0.35 1.515 0.44 ;
      RECT 0.56 0.95 0.749 1.04 ;
      RECT 0.659 0.645 0.749 1.04 ;
      RECT 0.659 0.645 0.845 0.735 ;
      RECT 0.755 0.35 0.845 0.735 ;
      RECT 0.66 0.35 0.845 0.44 ;
  END
END LATHRX1H7R

MACRO LATHRX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATHRX2H7R 0 0 ;
  SIZE 4.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.6 1.48 ;
        RECT 4.2 0.845 4.29 1.48 ;
        RECT 3.62 1.165 3.76 1.48 ;
        RECT 3.035 1.165 3.175 1.48 ;
        RECT 2.565 1.055 2.655 1.48 ;
        RECT 1.82 1.24 1.96 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.6 0.08 ;
        RECT 4.27 -0.08 4.36 0.34 ;
        RECT 3.75 -0.08 3.84 0.33 ;
        RECT 3.25 -0.08 3.34 0.33 ;
        RECT 2.02 -0.08 2.16 0.16 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.655 0.562 1.745 0.777 ;
        RECT 1.57 0.562 1.745 0.652 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.455 0.375 0.635 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END G
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.455 0.225 3.615 0.315 ;
        RECT 3.355 0.805 3.545 0.895 ;
        RECT 3.455 0.225 3.545 0.895 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.02 0.225 4.145 0.375 ;
        RECT 3.925 0.805 4.11 0.895 ;
        RECT 4.02 0.225 4.11 0.895 ;
        RECT 3.995 0.225 4.145 0.315 ;
      LAYER MET2 ;
        RECT 4.05 0.18 4.15 0.56 ;
      LAYER VIA1 ;
        RECT 4.055 0.255 4.145 0.345 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.96 0.455 2.175 0.545 ;
        RECT 1.96 0.455 2.05 0.63 ;
      LAYER MET2 ;
        RECT 2.05 0.23 2.15 0.76 ;
      LAYER VIA1 ;
        RECT 2.055 0.455 2.145 0.545 ;
    END
  END RN
  OBS
    LAYER MET1 ;
      RECT 3.055 0.985 3.725 1.075 ;
      RECT 3.635 0.535 3.725 1.075 ;
      RECT 3.055 0.295 3.145 1.075 ;
      RECT 2.365 0.82 3.145 0.91 ;
      RECT 3.635 0.535 3.93 0.627 ;
      RECT 3.84 0.487 3.93 0.627 ;
      RECT 3 0.295 3.145 0.435 ;
      RECT 1.089 0.96 1.623 1.05 ;
      RECT 1.089 0.96 1.709 0.987 ;
      RECT 1.089 0.96 1.713 0.962 ;
      RECT 2.185 0.64 2.275 0.96 ;
      RECT 1.663 0.87 2.275 0.96 ;
      RECT 1.573 0.937 2.275 0.96 ;
      RECT 1.623 0.89 1.663 1.03 ;
      RECT 1.089 0.35 1.179 1.05 ;
      RECT 1.619 0.912 2.275 0.96 ;
      RECT 2.185 0.64 2.965 0.73 ;
      RECT 2.82 0.57 2.965 0.73 ;
      RECT 2.82 0.25 2.91 0.73 ;
      RECT 0.965 0.35 1.179 0.44 ;
      RECT 2.72 0.25 2.91 0.34 ;
      RECT 0.045 0.725 0.16 1.065 ;
      RECT 0.045 0.725 0.569 0.815 ;
      RECT 0.479 0.675 0.569 0.815 ;
      RECT 0.045 0.275 0.135 1.065 ;
      RECT 2.507 0.46 2.73 0.55 ;
      RECT 2.507 0.25 2.597 0.55 ;
      RECT 0.045 0.275 0.517 0.365 ;
      RECT 1.748 0.25 2.597 0.34 ;
      RECT 1.707 0.19 1.748 0.32 ;
      RECT 1.668 0.25 2.597 0.28 ;
      RECT 0.479 0.256 0.622 0.279 ;
      RECT 0.563 0.18 0.584 0.309 ;
      RECT 0.584 0.17 1.707 0.26 ;
      RECT 0.517 0.214 0.563 0.342 ;
      RECT 0.517 0.23 1.787 0.26 ;
      RECT 2.205 1.06 2.295 1.23 ;
      RECT 0.839 1.14 1.699 1.23 ;
      RECT 0.839 1.14 1.779 1.169 ;
      RECT 1.741 1.06 2.295 1.15 ;
      RECT 1.661 1.121 2.295 1.15 ;
      RECT 1.699 1.081 1.741 1.209 ;
      RECT 0.839 0.847 0.929 1.23 ;
      RECT 1.375 0.78 1.534 0.87 ;
      RECT 1.375 0.35 1.465 0.87 ;
      RECT 1.375 0.35 1.515 0.44 ;
      RECT 0.56 0.905 0.749 0.995 ;
      RECT 0.659 0.645 0.749 0.995 ;
      RECT 0.659 0.645 0.845 0.735 ;
      RECT 0.755 0.35 0.845 0.735 ;
      RECT 0.705 0.35 0.845 0.44 ;
  END
END LATHRX2H7R

MACRO LATHSRX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATHSRX0P5H7R 0 0 ;
  SIZE 5.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.2 1.48 ;
        RECT 4.455 1.07 4.545 1.48 ;
        RECT 3.5 1.225 3.64 1.48 ;
        RECT 2.98 1.225 3.12 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.2 0.08 ;
        RECT 4.6 -0.08 4.74 0.175 ;
        RECT 3.68 -0.08 3.82 0.175 ;
        RECT 2.74 -0.08 2.88 0.175 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.425 0.425 1.545 0.65 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.55 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END G
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.255 0.36 4.395 0.45 ;
        RECT 4.255 0.36 4.345 0.601 ;
        RECT 4.146 0.628 4.255 0.679 ;
        RECT 4.19 0.583 4.301 0.646 ;
        RECT 4.236 0.55 4.255 0.679 ;
        RECT 4.1 0.673 4.236 0.711 ;
        RECT 4.1 0.673 4.19 0.945 ;
      LAYER MET2 ;
        RECT 4.25 0.225 4.35 0.76 ;
      LAYER VIA1 ;
        RECT 4.255 0.455 4.345 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.023 0.36 4.165 0.45 ;
        RECT 3.941 0.42 4.061 0.469 ;
        RECT 3.985 0.379 4.023 0.507 ;
        RECT 3.815 0.855 3.985 0.945 ;
        RECT 3.895 0.465 3.985 0.945 ;
      LAYER MET2 ;
        RECT 3.85 0.63 3.95 1.16 ;
      LAYER VIA1 ;
        RECT 3.855 0.855 3.945 0.945 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.61 0.605 2.76 0.785 ;
      LAYER MET2 ;
        RECT 2.65 0.43 2.75 0.96 ;
      LAYER VIA1 ;
        RECT 2.655 0.655 2.745 0.745 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.39 0.675 3.575 0.815 ;
        RECT 3.425 0.655 3.575 0.815 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 4.68 0.95 4.945 1.04 ;
      RECT 4.855 0.28 4.945 1.04 ;
      RECT 3.71 0.325 3.8 0.735 ;
      RECT 2.37 0.425 2.46 0.59 ;
      RECT 2.37 0.425 2.758 0.515 ;
      RECT 3.699 0.325 3.801 0.415 ;
      RECT 4.574 0.28 5.005 0.37 ;
      RECT 3.994 0.17 4.426 0.26 ;
      RECT 3.051 0.17 3.506 0.26 ;
      RECT 4.536 0.261 4.574 0.37 ;
      RECT 4.51 0.229 4.536 0.357 ;
      RECT 4.464 0.193 4.51 0.321 ;
      RECT 4.426 0.17 4.464 0.279 ;
      RECT 3.956 0.17 3.994 0.279 ;
      RECT 3.931 0.182 3.956 0.311 ;
      RECT 3.885 0.218 3.931 0.346 ;
      RECT 3.839 0.264 3.885 0.392 ;
      RECT 3.801 0.306 3.839 0.415 ;
      RECT 3.661 0.306 3.699 0.415 ;
      RECT 3.636 0.274 3.661 0.403 ;
      RECT 3.59 0.239 3.636 0.367 ;
      RECT 3.544 0.193 3.59 0.321 ;
      RECT 3.506 0.17 3.544 0.279 ;
      RECT 3.013 0.17 3.051 0.279 ;
      RECT 2.98 0.186 3.013 0.315 ;
      RECT 2.934 0.226 2.98 0.354 ;
      RECT 2.888 0.272 2.934 0.4 ;
      RECT 2.842 0.318 2.888 0.446 ;
      RECT 2.796 0.364 2.842 0.492 ;
      RECT 2.758 0.406 2.796 0.515 ;
      RECT 2.885 1.045 4.259 1.135 ;
      RECT 2.885 1.045 4.305 1.112 ;
      RECT 2.37 0.875 2.51 1.05 ;
      RECT 0.875 0.17 0.965 1.05 ;
      RECT 4.221 1.026 4.351 1.066 ;
      RECT 2.885 0.533 2.975 1.135 ;
      RECT 4.259 0.984 4.351 1.066 ;
      RECT 4.305 0.938 4.397 1.02 ;
      RECT 2.37 0.875 2.975 0.965 ;
      RECT 4.351 0.892 4.471 0.946 ;
      RECT 4.397 0.855 4.425 0.983 ;
      RECT 4.425 0.625 4.515 0.901 ;
      RECT 2.37 0.685 2.46 1.05 ;
      RECT 2.05 0.685 2.46 0.775 ;
      RECT 4.425 0.625 4.765 0.715 ;
      RECT 2.05 0.35 2.14 0.775 ;
      RECT 2.931 0.488 3.021 0.571 ;
      RECT 2.931 0.488 3.067 0.525 ;
      RECT 2.975 0.443 3.091 0.49 ;
      RECT 3.021 0.397 3.129 0.459 ;
      RECT 3.067 0.362 3.091 0.49 ;
      RECT 3.091 0.35 3.235 0.44 ;
      RECT 1.691 0.35 2.14 0.44 ;
      RECT 1.687 0.31 1.691 0.438 ;
      RECT 1.641 0.285 1.687 0.413 ;
      RECT 1.595 0.239 1.641 0.367 ;
      RECT 1.595 0.331 1.729 0.367 ;
      RECT 1.549 0.193 1.595 0.321 ;
      RECT 1.511 0.239 1.641 0.279 ;
      RECT 0.875 0.17 1.549 0.26 ;
      RECT 3.15 0.865 3.29 0.955 ;
      RECT 3.15 0.553 3.24 0.955 ;
      RECT 3.065 0.655 3.24 0.745 ;
      RECT 3.15 0.553 3.314 0.62 ;
      RECT 3.196 0.53 3.371 0.586 ;
      RECT 3.314 0.486 3.325 0.615 ;
      RECT 3.325 0.35 3.415 0.541 ;
      RECT 3.276 0.511 3.415 0.541 ;
      RECT 3.325 0.35 3.465 0.44 ;
      RECT 1.735 1.14 2.75 1.23 ;
      RECT 2.66 1.07 2.75 1.23 ;
      RECT 2.475 0.17 2.615 0.325 ;
      RECT 1.77 0.17 2.615 0.26 ;
      RECT 0.695 1.14 1.61 1.23 ;
      RECT 1.52 0.96 1.61 1.23 ;
      RECT 0.695 0.26 0.785 1.23 ;
      RECT 0.545 1.045 0.785 1.135 ;
      RECT 1.52 0.96 2.28 1.05 ;
      RECT 2.19 0.87 2.28 1.05 ;
      RECT 0.545 0.26 0.785 0.35 ;
      RECT 1.235 0.78 1.86 0.87 ;
      RECT 1.235 0.73 1.325 0.87 ;
      RECT 1.055 0.96 1.24 1.05 ;
      RECT 1.055 0.35 1.145 1.05 ;
      RECT 1.055 0.35 1.27 0.44 ;
      RECT 0.045 0.865 0.16 1.065 ;
      RECT 0.045 0.865 0.56 0.955 ;
      RECT 0.47 0.655 0.56 0.955 ;
      RECT 0.045 0.28 0.135 1.065 ;
      RECT 0.045 0.28 0.185 0.37 ;
  END
END LATHSRX0P5H7R

MACRO LATHSRX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATHSRX1H7R 0 0 ;
  SIZE 5.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.2 1.48 ;
        RECT 4.455 1.07 4.545 1.48 ;
        RECT 3.5 1.225 3.64 1.48 ;
        RECT 2.98 1.225 3.12 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.2 0.08 ;
        RECT 4.6 -0.08 4.74 0.175 ;
        RECT 3.68 -0.08 3.82 0.175 ;
        RECT 2.74 -0.08 2.88 0.175 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.425 0.425 1.545 0.65 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.55 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END G
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.255 0.36 4.395 0.45 ;
        RECT 4.255 0.36 4.345 0.601 ;
        RECT 4.146 0.628 4.255 0.679 ;
        RECT 4.19 0.583 4.301 0.646 ;
        RECT 4.236 0.55 4.255 0.679 ;
        RECT 4.1 0.673 4.236 0.711 ;
        RECT 4.1 0.673 4.19 0.945 ;
      LAYER MET2 ;
        RECT 4.25 0.225 4.35 0.76 ;
      LAYER VIA1 ;
        RECT 4.255 0.455 4.345 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.023 0.36 4.165 0.45 ;
        RECT 3.941 0.42 4.061 0.469 ;
        RECT 3.985 0.379 4.023 0.507 ;
        RECT 3.815 0.855 3.985 0.945 ;
        RECT 3.895 0.465 3.985 0.945 ;
      LAYER MET2 ;
        RECT 3.85 0.63 3.95 1.16 ;
      LAYER VIA1 ;
        RECT 3.855 0.855 3.945 0.945 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.61 0.605 2.76 0.785 ;
      LAYER MET2 ;
        RECT 2.65 0.43 2.75 0.96 ;
      LAYER VIA1 ;
        RECT 2.655 0.655 2.745 0.745 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.39 0.675 3.575 0.815 ;
        RECT 3.425 0.655 3.575 0.815 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 4.68 0.95 4.945 1.04 ;
      RECT 4.855 0.28 4.945 1.04 ;
      RECT 3.71 0.325 3.8 0.735 ;
      RECT 2.37 0.425 2.46 0.59 ;
      RECT 2.37 0.425 2.758 0.515 ;
      RECT 3.699 0.325 3.801 0.415 ;
      RECT 4.574 0.28 5.005 0.37 ;
      RECT 3.994 0.17 4.426 0.26 ;
      RECT 3.051 0.17 3.506 0.26 ;
      RECT 4.536 0.261 4.574 0.37 ;
      RECT 4.51 0.229 4.536 0.357 ;
      RECT 4.464 0.193 4.51 0.321 ;
      RECT 4.426 0.17 4.464 0.279 ;
      RECT 3.956 0.17 3.994 0.279 ;
      RECT 3.931 0.182 3.956 0.311 ;
      RECT 3.885 0.218 3.931 0.346 ;
      RECT 3.839 0.264 3.885 0.392 ;
      RECT 3.801 0.306 3.839 0.415 ;
      RECT 3.661 0.306 3.699 0.415 ;
      RECT 3.636 0.274 3.661 0.403 ;
      RECT 3.59 0.239 3.636 0.367 ;
      RECT 3.544 0.193 3.59 0.321 ;
      RECT 3.506 0.17 3.544 0.279 ;
      RECT 3.013 0.17 3.051 0.279 ;
      RECT 2.98 0.186 3.013 0.315 ;
      RECT 2.934 0.226 2.98 0.354 ;
      RECT 2.888 0.272 2.934 0.4 ;
      RECT 2.842 0.318 2.888 0.446 ;
      RECT 2.796 0.364 2.842 0.492 ;
      RECT 2.758 0.406 2.796 0.515 ;
      RECT 2.885 1.045 4.259 1.135 ;
      RECT 2.885 1.045 4.305 1.112 ;
      RECT 2.37 0.875 2.51 1.05 ;
      RECT 0.875 0.17 0.965 1.05 ;
      RECT 4.221 1.026 4.351 1.066 ;
      RECT 2.885 0.533 2.975 1.135 ;
      RECT 4.259 0.984 4.351 1.066 ;
      RECT 4.305 0.938 4.397 1.02 ;
      RECT 2.37 0.875 2.975 0.965 ;
      RECT 4.351 0.892 4.471 0.946 ;
      RECT 4.397 0.855 4.425 0.983 ;
      RECT 4.425 0.625 4.515 0.901 ;
      RECT 2.37 0.685 2.46 1.05 ;
      RECT 2.05 0.685 2.46 0.775 ;
      RECT 4.425 0.625 4.765 0.715 ;
      RECT 2.05 0.35 2.14 0.775 ;
      RECT 2.931 0.488 3.021 0.571 ;
      RECT 2.931 0.488 3.067 0.525 ;
      RECT 2.975 0.443 3.091 0.49 ;
      RECT 3.021 0.397 3.129 0.459 ;
      RECT 3.067 0.362 3.091 0.49 ;
      RECT 3.091 0.35 3.235 0.44 ;
      RECT 1.691 0.35 2.14 0.44 ;
      RECT 1.687 0.31 1.691 0.438 ;
      RECT 1.641 0.285 1.687 0.413 ;
      RECT 1.595 0.239 1.641 0.367 ;
      RECT 1.595 0.331 1.729 0.367 ;
      RECT 1.549 0.193 1.595 0.321 ;
      RECT 1.511 0.239 1.641 0.279 ;
      RECT 0.875 0.17 1.549 0.26 ;
      RECT 3.15 0.865 3.29 0.955 ;
      RECT 3.15 0.553 3.24 0.955 ;
      RECT 3.065 0.655 3.24 0.745 ;
      RECT 3.15 0.553 3.314 0.62 ;
      RECT 3.196 0.53 3.371 0.586 ;
      RECT 3.314 0.486 3.325 0.615 ;
      RECT 3.325 0.35 3.415 0.541 ;
      RECT 3.276 0.511 3.415 0.541 ;
      RECT 3.325 0.35 3.465 0.44 ;
      RECT 1.735 1.14 2.75 1.23 ;
      RECT 2.66 1.07 2.75 1.23 ;
      RECT 2.475 0.17 2.615 0.325 ;
      RECT 1.77 0.17 2.615 0.26 ;
      RECT 0.695 1.14 1.61 1.23 ;
      RECT 1.52 0.96 1.61 1.23 ;
      RECT 0.695 0.26 0.785 1.23 ;
      RECT 0.545 1.045 0.785 1.135 ;
      RECT 1.52 0.96 2.28 1.05 ;
      RECT 2.19 0.87 2.28 1.05 ;
      RECT 0.545 0.26 0.785 0.35 ;
      RECT 1.235 0.78 1.86 0.87 ;
      RECT 1.235 0.73 1.325 0.87 ;
      RECT 1.055 0.96 1.24 1.05 ;
      RECT 1.055 0.35 1.145 1.05 ;
      RECT 1.055 0.35 1.27 0.44 ;
      RECT 0.045 0.865 0.16 1.065 ;
      RECT 0.045 0.865 0.56 0.955 ;
      RECT 0.47 0.655 0.56 0.955 ;
      RECT 0.045 0.28 0.135 1.065 ;
      RECT 0.045 0.28 0.185 0.37 ;
  END
END LATHSRX1H7R

MACRO LATHSRX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATHSRX2H7R 0 0 ;
  SIZE 5.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.2 1.48 ;
        RECT 4.455 1.07 4.545 1.48 ;
        RECT 3.5 1.225 3.64 1.48 ;
        RECT 2.98 1.225 3.12 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.2 0.08 ;
        RECT 4.6 -0.08 4.74 0.175 ;
        RECT 3.68 -0.08 3.82 0.175 ;
        RECT 2.74 -0.08 2.88 0.175 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.425 0.425 1.545 0.65 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.55 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END G
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.255 0.36 4.395 0.45 ;
        RECT 4.255 0.36 4.345 0.601 ;
        RECT 4.146 0.628 4.255 0.679 ;
        RECT 4.19 0.583 4.301 0.646 ;
        RECT 4.236 0.55 4.255 0.679 ;
        RECT 4.1 0.673 4.236 0.711 ;
        RECT 4.1 0.673 4.19 0.945 ;
      LAYER MET2 ;
        RECT 4.25 0.225 4.35 0.76 ;
      LAYER VIA1 ;
        RECT 4.255 0.455 4.345 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.023 0.36 4.165 0.45 ;
        RECT 3.941 0.42 4.061 0.469 ;
        RECT 3.985 0.379 4.023 0.507 ;
        RECT 3.815 0.855 3.985 0.945 ;
        RECT 3.895 0.465 3.985 0.945 ;
      LAYER MET2 ;
        RECT 3.85 0.63 3.95 1.16 ;
      LAYER VIA1 ;
        RECT 3.855 0.855 3.945 0.945 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.61 0.605 2.76 0.785 ;
      LAYER MET2 ;
        RECT 2.65 0.43 2.75 0.96 ;
      LAYER VIA1 ;
        RECT 2.655 0.655 2.745 0.745 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.39 0.675 3.575 0.815 ;
        RECT 3.425 0.655 3.575 0.815 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 4.68 0.95 4.945 1.04 ;
      RECT 4.855 0.28 4.945 1.04 ;
      RECT 3.71 0.325 3.8 0.735 ;
      RECT 2.37 0.425 2.46 0.59 ;
      RECT 2.37 0.425 2.758 0.515 ;
      RECT 3.699 0.325 3.801 0.415 ;
      RECT 4.574 0.28 5.005 0.37 ;
      RECT 3.994 0.17 4.426 0.26 ;
      RECT 3.051 0.17 3.506 0.26 ;
      RECT 4.536 0.261 4.574 0.37 ;
      RECT 4.51 0.229 4.536 0.357 ;
      RECT 4.464 0.193 4.51 0.321 ;
      RECT 4.426 0.17 4.464 0.279 ;
      RECT 3.956 0.17 3.994 0.279 ;
      RECT 3.931 0.182 3.956 0.311 ;
      RECT 3.885 0.218 3.931 0.346 ;
      RECT 3.839 0.264 3.885 0.392 ;
      RECT 3.801 0.306 3.839 0.415 ;
      RECT 3.661 0.306 3.699 0.415 ;
      RECT 3.636 0.274 3.661 0.403 ;
      RECT 3.59 0.239 3.636 0.367 ;
      RECT 3.544 0.193 3.59 0.321 ;
      RECT 3.506 0.17 3.544 0.279 ;
      RECT 3.013 0.17 3.051 0.279 ;
      RECT 2.98 0.186 3.013 0.315 ;
      RECT 2.934 0.226 2.98 0.354 ;
      RECT 2.888 0.272 2.934 0.4 ;
      RECT 2.842 0.318 2.888 0.446 ;
      RECT 2.796 0.364 2.842 0.492 ;
      RECT 2.758 0.406 2.796 0.515 ;
      RECT 2.885 1.045 4.259 1.135 ;
      RECT 2.885 1.045 4.305 1.112 ;
      RECT 2.37 0.875 2.51 1.05 ;
      RECT 4.221 1.026 4.351 1.066 ;
      RECT 2.885 0.533 2.975 1.135 ;
      RECT 4.259 0.984 4.351 1.066 ;
      RECT 0.875 0.17 0.965 1.005 ;
      RECT 4.305 0.938 4.397 1.02 ;
      RECT 2.37 0.875 2.975 0.965 ;
      RECT 4.351 0.892 4.471 0.946 ;
      RECT 4.397 0.855 4.425 0.983 ;
      RECT 4.425 0.625 4.515 0.901 ;
      RECT 2.37 0.685 2.46 1.05 ;
      RECT 2.05 0.685 2.46 0.775 ;
      RECT 4.425 0.625 4.765 0.715 ;
      RECT 2.05 0.35 2.14 0.775 ;
      RECT 2.931 0.488 3.021 0.571 ;
      RECT 2.931 0.488 3.067 0.525 ;
      RECT 2.975 0.443 3.091 0.49 ;
      RECT 3.021 0.397 3.129 0.459 ;
      RECT 3.067 0.362 3.091 0.49 ;
      RECT 3.091 0.35 3.235 0.44 ;
      RECT 1.691 0.35 2.14 0.44 ;
      RECT 1.687 0.31 1.691 0.438 ;
      RECT 1.641 0.285 1.687 0.413 ;
      RECT 1.595 0.239 1.641 0.367 ;
      RECT 1.595 0.331 1.729 0.367 ;
      RECT 1.549 0.193 1.595 0.321 ;
      RECT 1.511 0.239 1.641 0.279 ;
      RECT 0.875 0.17 1.549 0.26 ;
      RECT 3.15 0.865 3.29 0.955 ;
      RECT 3.15 0.553 3.24 0.955 ;
      RECT 3.065 0.655 3.24 0.745 ;
      RECT 3.15 0.553 3.314 0.62 ;
      RECT 3.196 0.53 3.371 0.586 ;
      RECT 3.314 0.486 3.325 0.615 ;
      RECT 3.325 0.35 3.415 0.541 ;
      RECT 3.276 0.511 3.415 0.541 ;
      RECT 3.325 0.35 3.465 0.44 ;
      RECT 1.735 1.14 2.75 1.23 ;
      RECT 2.66 1.07 2.75 1.23 ;
      RECT 2.475 0.17 2.615 0.325 ;
      RECT 1.77 0.17 2.615 0.26 ;
      RECT 0.695 1.14 1.61 1.23 ;
      RECT 1.52 0.96 1.61 1.23 ;
      RECT 0.695 0.26 0.785 1.23 ;
      RECT 0.545 1.045 0.785 1.135 ;
      RECT 1.52 0.96 2.28 1.05 ;
      RECT 2.19 0.87 2.28 1.05 ;
      RECT 0.545 0.26 0.785 0.35 ;
      RECT 1.235 0.78 1.86 0.87 ;
      RECT 1.235 0.73 1.325 0.87 ;
      RECT 1.055 0.96 1.24 1.05 ;
      RECT 1.055 0.35 1.145 1.05 ;
      RECT 1.055 0.35 1.24 0.44 ;
      RECT 0.045 0.865 0.16 1.065 ;
      RECT 0.045 0.865 0.56 0.955 ;
      RECT 0.47 0.655 0.56 0.955 ;
      RECT 0.045 0.28 0.135 1.065 ;
      RECT 0.045 0.28 0.185 0.37 ;
  END
END LATHSRX2H7R

MACRO LATHSX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATHSX0P5H7R 0 0 ;
  SIZE 5.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.4 1.48 ;
        RECT 4.89 1.05 4.98 1.48 ;
        RECT 3.939 1.2 4.029 1.48 ;
        RECT 2.555 1.113 2.695 1.48 ;
        RECT 0.802 1.225 0.942 1.48 ;
        RECT 0.32 1.015 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.4 0.08 ;
        RECT 4.886 -0.08 5.026 0.175 ;
        RECT 3.655 -0.08 3.745 0.33 ;
        RECT 2.425 -0.08 2.565 0.36 ;
        RECT 0.8 -0.08 0.89 0.33 ;
        RECT 0.32 -0.08 0.41 0.345 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.147 0.68 1.287 0.77 ;
        RECT 1.147 0.455 1.237 0.77 ;
        RECT 0.705 0.455 1.237 0.555 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.565 0.425 3.745 0.575 ;
      LAYER MET2 ;
        RECT 3.65 0.23 3.75 0.76 ;
      LAYER VIA1 ;
        RECT 3.655 0.455 3.745 0.545 ;
    END
  END G
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.64 0.87 4.93 0.96 ;
        RECT 4.84 0.455 4.93 0.96 ;
        RECT 4.535 0.455 4.93 0.545 ;
        RECT 4.64 0.87 4.73 1.045 ;
        RECT 4.535 0.35 4.675 0.545 ;
      LAYER MET2 ;
        RECT 4.65 0.225 4.75 0.76 ;
      LAYER VIA1 ;
        RECT 4.655 0.455 4.745 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.219 0.504 4.345 0.92 ;
        RECT 4.219 0.464 4.311 0.92 ;
        RECT 4.174 0.418 4.265 0.5 ;
        RECT 4.034 0.372 4.219 0.44 ;
        RECT 4.034 0.35 4.174 0.44 ;
        RECT 4.136 0.418 4.265 0.459 ;
      LAYER MET2 ;
        RECT 4.25 0.425 4.35 0.96 ;
      LAYER VIA1 ;
        RECT 4.255 0.655 4.345 0.745 ;
    END
  END QN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.455 0.375 0.635 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 3.022 0.96 3.695 1.05 ;
      RECT 5.176 0.265 5.266 1.045 ;
      RECT 2.994 0.908 3.022 1.036 ;
      RECT 2.994 0.96 3.741 1.027 ;
      RECT 2.948 0.871 2.994 0.999 ;
      RECT 3.653 0.939 3.787 0.981 ;
      RECT 2.948 0.941 3.06 0.999 ;
      RECT 2.902 0.825 2.948 0.953 ;
      RECT 3.695 0.895 3.787 0.981 ;
      RECT 3.695 0.895 3.833 0.935 ;
      RECT 2.856 0.779 2.902 0.907 ;
      RECT 3.741 0.849 3.854 0.902 ;
      RECT 2.81 0.733 2.856 0.861 ;
      RECT 3.787 0.803 3.9 0.868 ;
      RECT 3.833 0.769 3.854 0.902 ;
      RECT 3.854 0.17 3.944 0.823 ;
      RECT 2.772 0.779 2.902 0.819 ;
      RECT 2.13 0.71 2.81 0.8 ;
      RECT 3.854 0.576 4.034 0.666 ;
      RECT 4.81 0.265 5.266 0.355 ;
      RECT 4.799 0.221 4.81 0.35 ;
      RECT 4.753 0.193 4.799 0.321 ;
      RECT 4.715 0.246 4.848 0.279 ;
      RECT 3.854 0.17 4.753 0.26 ;
      RECT 2.785 1.14 3.779 1.23 ;
      RECT 2.785 1.14 3.825 1.207 ;
      RECT 3.737 1.119 3.867 1.163 ;
      RECT 2.785 1.013 2.875 1.23 ;
      RECT 3.779 1.075 3.909 1.121 ;
      RECT 3.825 1.031 3.867 1.163 ;
      RECT 4.435 0.635 4.525 1.1 ;
      RECT 3.867 1.01 4.525 1.1 ;
      RECT 2.776 0.94 2.785 1.069 ;
      RECT 2.73 0.913 2.776 1.041 ;
      RECT 2.73 0.968 2.831 1.041 ;
      RECT 2.692 0.968 2.831 0.999 ;
      RECT 1.56 0.89 2.73 0.98 ;
      RECT 1.56 0.53 1.65 0.98 ;
      RECT 4.435 0.635 4.75 0.725 ;
      RECT 1.56 0.53 1.857 0.62 ;
      RECT 1.767 0.17 1.857 0.62 ;
      RECT 1.767 0.17 1.897 0.365 ;
      RECT 1.121 0.17 1.261 0.305 ;
      RECT 1.121 0.17 1.897 0.26 ;
      RECT 3.47 0.78 3.612 0.87 ;
      RECT 3.467 0.696 3.47 0.825 ;
      RECT 3.421 0.672 3.467 0.8 ;
      RECT 3.421 0.762 3.552 0.8 ;
      RECT 3.421 0.721 3.516 0.8 ;
      RECT 3.375 0.626 3.421 0.754 ;
      RECT 3.329 0.58 3.375 0.708 ;
      RECT 3.285 0.171 3.329 0.663 ;
      RECT 3.239 0.171 3.329 0.618 ;
      RECT 2.868 0.171 3.329 0.261 ;
      RECT 3.1 0.78 3.255 0.87 ;
      RECT 3.066 0.725 3.1 0.853 ;
      RECT 3.02 0.685 3.066 0.813 ;
      RECT 1.742 0.71 2.04 0.8 ;
      RECT 1.95 0.45 2.04 0.8 ;
      RECT 3.02 0.761 3.138 0.813 ;
      RECT 2.974 0.639 3.02 0.767 ;
      RECT 2.928 0.593 2.974 0.721 ;
      RECT 2.882 0.547 2.928 0.675 ;
      RECT 2.836 0.501 2.882 0.629 ;
      RECT 2.79 0.455 2.836 0.583 ;
      RECT 2.77 0.31 2.79 0.55 ;
      RECT 2.7 0.31 2.79 0.54 ;
      RECT 1.95 0.45 2.79 0.54 ;
      RECT 1.065 1.07 2.448 1.16 ;
      RECT 0.532 1.045 0.672 1.15 ;
      RECT 0.532 1.045 1.155 1.135 ;
      RECT 1.277 0.865 1.467 0.98 ;
      RECT 1.377 0.35 1.467 0.98 ;
      RECT 0.879 0.865 1.467 0.955 ;
      RECT 0.879 0.645 0.969 0.955 ;
      RECT 0.525 0.645 0.969 0.735 ;
      RECT 0.525 0.28 0.615 0.735 ;
      RECT 1.377 0.35 1.677 0.44 ;
      RECT 0.525 0.28 0.665 0.37 ;
      RECT 0.045 0.825 0.16 1.025 ;
      RECT 0.045 0.825 0.777 0.915 ;
      RECT 0.045 0.28 0.135 1.025 ;
      RECT 0.045 0.28 0.185 0.37 ;
  END
END LATHSX0P5H7R

MACRO LATHSX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATHSX1H7R 0 0 ;
  SIZE 5.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.4 1.48 ;
        RECT 4.89 1.05 4.98 1.48 ;
        RECT 3.939 1.2 4.029 1.48 ;
        RECT 2.555 1.113 2.695 1.48 ;
        RECT 0.802 1.225 0.942 1.48 ;
        RECT 0.32 1.015 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.4 0.08 ;
        RECT 4.886 -0.08 5.026 0.175 ;
        RECT 3.655 -0.08 3.745 0.33 ;
        RECT 2.425 -0.08 2.565 0.36 ;
        RECT 0.8 -0.08 0.89 0.33 ;
        RECT 0.32 -0.08 0.41 0.345 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.147 0.68 1.287 0.77 ;
        RECT 1.147 0.455 1.237 0.77 ;
        RECT 0.705 0.455 1.237 0.555 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.565 0.425 3.745 0.575 ;
      LAYER MET2 ;
        RECT 3.65 0.23 3.75 0.76 ;
      LAYER VIA1 ;
        RECT 3.655 0.455 3.745 0.545 ;
    END
  END G
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.615 0.87 4.93 0.96 ;
        RECT 4.84 0.455 4.93 0.96 ;
        RECT 4.535 0.455 4.93 0.545 ;
        RECT 4.535 0.35 4.675 0.545 ;
      LAYER MET2 ;
        RECT 4.65 0.225 4.75 0.76 ;
      LAYER VIA1 ;
        RECT 4.655 0.455 4.745 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.219 0.504 4.345 0.92 ;
        RECT 4.219 0.464 4.311 0.92 ;
        RECT 4.174 0.418 4.265 0.5 ;
        RECT 4.034 0.372 4.219 0.44 ;
        RECT 4.034 0.35 4.174 0.44 ;
        RECT 4.136 0.418 4.265 0.459 ;
      LAYER MET2 ;
        RECT 4.25 0.425 4.35 0.96 ;
      LAYER VIA1 ;
        RECT 4.255 0.655 4.345 0.745 ;
    END
  END QN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.455 0.375 0.635 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 3.022 0.96 3.695 1.05 ;
      RECT 5.176 0.265 5.266 1.045 ;
      RECT 2.994 0.908 3.022 1.036 ;
      RECT 2.994 0.96 3.741 1.027 ;
      RECT 2.948 0.871 2.994 0.999 ;
      RECT 3.653 0.939 3.787 0.981 ;
      RECT 2.948 0.941 3.06 0.999 ;
      RECT 2.902 0.825 2.948 0.953 ;
      RECT 3.695 0.895 3.787 0.981 ;
      RECT 3.695 0.895 3.833 0.935 ;
      RECT 2.856 0.779 2.902 0.907 ;
      RECT 3.741 0.849 3.854 0.902 ;
      RECT 2.81 0.733 2.856 0.861 ;
      RECT 3.787 0.803 3.9 0.868 ;
      RECT 3.833 0.769 3.854 0.902 ;
      RECT 3.854 0.17 3.944 0.823 ;
      RECT 2.772 0.779 2.902 0.819 ;
      RECT 2.13 0.71 2.81 0.8 ;
      RECT 3.854 0.576 4.034 0.666 ;
      RECT 4.81 0.265 5.266 0.355 ;
      RECT 4.799 0.221 4.81 0.35 ;
      RECT 4.753 0.193 4.799 0.321 ;
      RECT 4.715 0.246 4.848 0.279 ;
      RECT 3.854 0.17 4.753 0.26 ;
      RECT 2.785 1.14 3.779 1.23 ;
      RECT 2.785 1.14 3.825 1.207 ;
      RECT 3.737 1.119 3.867 1.163 ;
      RECT 2.785 1.013 2.875 1.23 ;
      RECT 3.779 1.075 3.909 1.121 ;
      RECT 3.825 1.031 3.867 1.163 ;
      RECT 4.435 0.635 4.525 1.1 ;
      RECT 3.867 1.01 4.525 1.1 ;
      RECT 2.776 0.94 2.785 1.069 ;
      RECT 2.73 0.913 2.776 1.041 ;
      RECT 2.73 0.968 2.831 1.041 ;
      RECT 2.692 0.968 2.831 0.999 ;
      RECT 1.56 0.89 2.73 0.98 ;
      RECT 1.56 0.53 1.65 0.98 ;
      RECT 4.435 0.635 4.75 0.725 ;
      RECT 1.56 0.53 1.857 0.62 ;
      RECT 1.767 0.17 1.857 0.62 ;
      RECT 1.767 0.17 1.897 0.365 ;
      RECT 1.121 0.17 1.261 0.305 ;
      RECT 1.121 0.17 1.897 0.26 ;
      RECT 3.47 0.78 3.612 0.87 ;
      RECT 3.467 0.696 3.47 0.825 ;
      RECT 3.421 0.672 3.467 0.8 ;
      RECT 3.421 0.762 3.552 0.8 ;
      RECT 3.421 0.721 3.516 0.8 ;
      RECT 3.375 0.626 3.421 0.754 ;
      RECT 3.329 0.58 3.375 0.708 ;
      RECT 3.285 0.171 3.329 0.663 ;
      RECT 3.239 0.171 3.329 0.618 ;
      RECT 2.868 0.171 3.329 0.261 ;
      RECT 3.1 0.78 3.255 0.87 ;
      RECT 3.066 0.725 3.1 0.853 ;
      RECT 3.02 0.685 3.066 0.813 ;
      RECT 1.742 0.71 2.04 0.8 ;
      RECT 1.95 0.45 2.04 0.8 ;
      RECT 3.02 0.761 3.138 0.813 ;
      RECT 2.974 0.639 3.02 0.767 ;
      RECT 2.928 0.593 2.974 0.721 ;
      RECT 2.882 0.547 2.928 0.675 ;
      RECT 2.836 0.501 2.882 0.629 ;
      RECT 2.79 0.455 2.836 0.583 ;
      RECT 2.77 0.31 2.79 0.55 ;
      RECT 2.7 0.31 2.79 0.54 ;
      RECT 1.95 0.45 2.79 0.54 ;
      RECT 1.065 1.07 2.448 1.16 ;
      RECT 0.532 1.045 0.672 1.15 ;
      RECT 0.532 1.045 1.155 1.135 ;
      RECT 1.277 0.865 1.467 0.98 ;
      RECT 1.377 0.35 1.467 0.98 ;
      RECT 0.879 0.865 1.467 0.955 ;
      RECT 0.879 0.645 0.969 0.955 ;
      RECT 0.525 0.645 0.969 0.735 ;
      RECT 0.525 0.28 0.615 0.735 ;
      RECT 1.377 0.35 1.677 0.44 ;
      RECT 0.525 0.28 0.665 0.37 ;
      RECT 0.045 0.825 0.16 1.025 ;
      RECT 0.045 0.825 0.777 0.915 ;
      RECT 0.045 0.28 0.135 1.025 ;
      RECT 0.045 0.28 0.185 0.37 ;
  END
END LATHSX1H7R

MACRO LATHSX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATHSX2H7R 0 0 ;
  SIZE 5.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.6 1.48 ;
        RECT 5.1 1.05 5.19 1.48 ;
        RECT 4.474 1.19 4.614 1.48 ;
        RECT 3.939 1.2 4.029 1.48 ;
        RECT 2.555 1.113 2.695 1.48 ;
        RECT 0.802 1.225 0.942 1.48 ;
        RECT 0.32 1.015 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.6 0.08 ;
        RECT 5.12 -0.08 5.26 0.175 ;
        RECT 4.389 -0.08 4.529 0.16 ;
        RECT 3.655 -0.08 3.745 0.33 ;
        RECT 2.425 -0.08 2.565 0.35 ;
        RECT 0.8 -0.08 0.89 0.33 ;
        RECT 0.32 -0.08 0.41 0.345 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.147 0.68 1.287 0.77 ;
        RECT 1.147 0.455 1.237 0.77 ;
        RECT 0.705 0.455 1.237 0.555 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.565 0.425 3.745 0.575 ;
      LAYER MET2 ;
        RECT 3.65 0.23 3.75 0.76 ;
      LAYER VIA1 ;
        RECT 3.655 0.455 3.745 0.545 ;
    END
  END G
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.85 0.87 5.2 0.96 ;
        RECT 5.11 0.455 5.2 0.96 ;
        RECT 4.769 0.455 5.2 0.545 ;
        RECT 4.85 0.87 4.94 1.11 ;
        RECT 4.769 0.35 4.909 0.545 ;
      LAYER MET2 ;
        RECT 4.85 0.23 4.95 0.76 ;
      LAYER VIA1 ;
        RECT 4.855 0.455 4.945 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.219 0.504 4.345 0.92 ;
        RECT 4.219 0.464 4.311 0.92 ;
        RECT 4.174 0.418 4.265 0.5 ;
        RECT 4.034 0.372 4.219 0.44 ;
        RECT 4.034 0.35 4.174 0.44 ;
        RECT 4.136 0.418 4.265 0.459 ;
      LAYER MET2 ;
        RECT 4.25 0.425 4.35 0.96 ;
      LAYER VIA1 ;
        RECT 4.255 0.655 4.345 0.745 ;
    END
  END QN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.455 0.375 0.635 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 3.06 0.96 3.653 1.05 ;
      RECT 5.41 0.265 5.5 1.045 ;
      RECT 2.13 0.71 2.772 0.8 ;
      RECT 3.944 0.576 4.034 0.666 ;
      RECT 5.082 0.265 5.5 0.355 ;
      RECT 4.347 0.25 4.611 0.34 ;
      RECT 4.731 0.17 4.949 0.26 ;
      RECT 3.944 0.17 4.212 0.26 ;
      RECT 5.044 0.246 5.082 0.355 ;
      RECT 5.033 0.221 5.044 0.35 ;
      RECT 4.987 0.193 5.033 0.321 ;
      RECT 4.949 0.17 4.987 0.279 ;
      RECT 4.691 0.17 4.731 0.28 ;
      RECT 4.651 0.19 4.691 0.32 ;
      RECT 4.611 0.23 4.651 0.34 ;
      RECT 4.338 0.245 4.347 0.34 ;
      RECT 4.292 0.218 4.338 0.34 ;
      RECT 4.267 0.182 4.292 0.328 ;
      RECT 4.258 0.17 4.267 0.311 ;
      RECT 4.212 0.17 4.258 0.283 ;
      RECT 3.9 0.17 3.944 0.823 ;
      RECT 3.854 0.17 3.9 0.868 ;
      RECT 3.833 0.769 3.854 0.902 ;
      RECT 3.787 0.803 3.833 0.935 ;
      RECT 3.741 0.849 3.787 0.981 ;
      RECT 3.695 0.895 3.741 1.027 ;
      RECT 3.653 0.939 3.695 1.05 ;
      RECT 3.022 0.941 3.06 1.05 ;
      RECT 2.994 0.908 3.022 1.036 ;
      RECT 2.948 0.871 2.994 0.999 ;
      RECT 2.902 0.825 2.948 0.953 ;
      RECT 2.856 0.779 2.902 0.907 ;
      RECT 2.81 0.733 2.856 0.861 ;
      RECT 2.772 0.71 2.81 0.819 ;
      RECT 2.785 1.14 3.779 1.23 ;
      RECT 2.785 1.14 3.825 1.207 ;
      RECT 3.737 1.119 3.867 1.163 ;
      RECT 2.785 1.013 2.875 1.23 ;
      RECT 3.779 1.075 3.909 1.121 ;
      RECT 3.825 1.031 3.867 1.163 ;
      RECT 4.669 0.69 4.759 1.1 ;
      RECT 3.867 1.01 4.759 1.1 ;
      RECT 2.776 0.94 2.785 1.069 ;
      RECT 2.73 0.913 2.776 1.041 ;
      RECT 2.73 0.968 2.831 1.041 ;
      RECT 2.692 0.968 2.831 0.999 ;
      RECT 1.56 0.89 2.73 0.98 ;
      RECT 1.56 0.53 1.65 0.98 ;
      RECT 4.669 0.69 5.019 0.78 ;
      RECT 1.56 0.53 1.857 0.62 ;
      RECT 1.767 0.17 1.857 0.62 ;
      RECT 1.767 0.17 1.897 0.365 ;
      RECT 1.121 0.17 1.261 0.305 ;
      RECT 1.121 0.17 1.897 0.26 ;
      RECT 3.47 0.78 3.612 0.87 ;
      RECT 3.467 0.696 3.47 0.825 ;
      RECT 3.421 0.672 3.467 0.8 ;
      RECT 3.421 0.762 3.552 0.8 ;
      RECT 3.421 0.721 3.516 0.8 ;
      RECT 3.375 0.626 3.421 0.754 ;
      RECT 3.329 0.58 3.375 0.708 ;
      RECT 3.285 0.171 3.329 0.663 ;
      RECT 3.239 0.171 3.329 0.618 ;
      RECT 2.863 0.171 3.329 0.261 ;
      RECT 3.13 0.78 3.285 0.87 ;
      RECT 3.091 0.722 3.13 0.851 ;
      RECT 3.045 0.68 3.091 0.808 ;
      RECT 1.742 0.71 2.04 0.8 ;
      RECT 1.95 0.44 2.04 0.8 ;
      RECT 3.045 0.761 3.168 0.808 ;
      RECT 2.999 0.634 3.045 0.762 ;
      RECT 2.953 0.588 2.999 0.716 ;
      RECT 2.907 0.542 2.953 0.67 ;
      RECT 2.861 0.496 2.907 0.624 ;
      RECT 2.815 0.45 2.861 0.578 ;
      RECT 2.79 0.35 2.815 0.543 ;
      RECT 2.675 0.35 2.815 0.53 ;
      RECT 1.95 0.44 2.815 0.53 ;
      RECT 1.065 1.07 2.448 1.16 ;
      RECT 0.532 1.045 0.672 1.15 ;
      RECT 0.532 1.045 1.155 1.135 ;
      RECT 1.277 0.865 1.467 0.98 ;
      RECT 1.377 0.35 1.467 0.98 ;
      RECT 0.879 0.865 1.467 0.955 ;
      RECT 0.879 0.645 0.969 0.955 ;
      RECT 0.525 0.645 0.969 0.735 ;
      RECT 0.525 0.28 0.615 0.735 ;
      RECT 1.377 0.35 1.677 0.44 ;
      RECT 0.525 0.28 0.665 0.37 ;
      RECT 0.045 0.825 0.16 1.025 ;
      RECT 0.045 0.825 0.777 0.915 ;
      RECT 0.045 0.28 0.135 1.025 ;
      RECT 0.045 0.28 0.185 0.37 ;
  END
END LATHSX2H7R

MACRO LATHX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATHX0P5H7R 0 0 ;
  SIZE 3.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.2 1.48 ;
        RECT 2.658 1.225 2.798 1.48 ;
        RECT 1.881 1.24 2.021 1.48 ;
        RECT 0.806 1.209 0.946 1.48 ;
        RECT 0.311 1.225 0.451 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.2 0.08 ;
        RECT 2.698 -0.08 2.788 0.362 ;
        RECT 1.851 -0.08 1.941 0.33 ;
        RECT 0.806 -0.08 0.946 0.204 ;
        RECT 0.32 -0.08 0.41 0.345 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.625 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.625 0.35 0.895 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END G
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.948 0.287 3.038 0.98 ;
        RECT 2.825 0.455 3.038 0.545 ;
      LAYER MET2 ;
        RECT 2.85 0.23 2.95 0.76 ;
      LAYER VIA1 ;
        RECT 2.855 0.455 2.945 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.055 0.872 2.302 0.962 ;
        RECT 2.055 0.28 2.241 0.37 ;
        RECT 2.055 0.28 2.145 0.962 ;
      LAYER MET2 ;
        RECT 2.05 0.23 2.15 0.76 ;
      LAYER VIA1 ;
        RECT 2.055 0.455 2.145 0.545 ;
    END
  END QN
  OBS
    LAYER MET1 ;
      RECT 1.287 1.059 2.598 1.149 ;
      RECT 1.287 1.059 2.644 1.126 ;
      RECT 2.56 1.04 2.673 1.089 ;
      RECT 1.819 0.687 1.909 1.149 ;
      RECT 2.598 0.998 2.719 1.051 ;
      RECT 2.644 0.96 2.673 1.089 ;
      RECT 2.673 0.63 2.763 1.006 ;
      RECT 1.671 0.687 1.909 0.777 ;
      RECT 1.671 0.241 1.761 0.777 ;
      RECT 1.318 0.241 1.761 0.331 ;
      RECT 2.392 0.285 2.532 0.955 ;
      RECT 2.307 0.598 2.532 0.738 ;
      RECT 1.491 0.879 1.631 0.969 ;
      RECT 0.541 0.84 0.796 0.93 ;
      RECT 0.706 0.294 0.796 0.93 ;
      RECT 1.491 0.445 1.581 0.969 ;
      RECT 1.222 0.445 1.581 0.555 ;
      RECT 0.706 0.445 1.581 0.535 ;
      RECT 0.541 0.294 0.796 0.384 ;
      RECT 0.07 1.02 1.085 1.11 ;
      RECT 0.07 1.02 1.131 1.087 ;
      RECT 1.047 1.001 1.177 1.041 ;
      RECT 0.07 0.255 0.16 1.11 ;
      RECT 1.085 0.959 1.177 1.041 ;
      RECT 1.131 0.913 1.223 0.995 ;
      RECT 1.177 0.867 1.297 0.921 ;
      RECT 1.223 0.83 1.251 0.958 ;
      RECT 1.251 0.67 1.341 0.876 ;
      RECT 0.526 0.569 0.616 0.745 ;
      RECT 0.516 0.496 0.526 0.624 ;
      RECT 0.47 0.468 0.516 0.596 ;
      RECT 0.47 0.524 0.572 0.596 ;
      RECT 0.432 0.524 0.572 0.554 ;
      RECT 0.07 0.445 0.47 0.535 ;
  END
END LATHX0P5H7R

MACRO LATHX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATHX1H7R 0 0 ;
  SIZE 3.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.2 1.48 ;
        RECT 2.658 1.225 2.798 1.48 ;
        RECT 1.881 1.24 2.021 1.48 ;
        RECT 0.806 1.209 0.946 1.48 ;
        RECT 0.311 1.225 0.451 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.2 0.08 ;
        RECT 2.698 -0.08 2.788 0.335 ;
        RECT 1.851 -0.08 1.941 0.35 ;
        RECT 0.806 -0.08 0.946 0.204 ;
        RECT 0.295 -0.08 0.435 0.352 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.625 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.625 0.35 0.895 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END G
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.948 0.287 3.038 0.98 ;
        RECT 2.825 0.455 3.038 0.545 ;
      LAYER MET2 ;
        RECT 2.85 0.23 2.95 0.76 ;
      LAYER VIA1 ;
        RECT 2.855 0.455 2.945 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.055 0.872 2.302 0.962 ;
        RECT 2.055 0.335 2.216 0.425 ;
        RECT 2.055 0.335 2.145 0.962 ;
      LAYER MET2 ;
        RECT 2.05 0.23 2.15 0.76 ;
      LAYER VIA1 ;
        RECT 2.055 0.455 2.145 0.545 ;
    END
  END QN
  OBS
    LAYER MET1 ;
      RECT 1.287 1.059 2.598 1.149 ;
      RECT 1.287 1.059 2.644 1.126 ;
      RECT 2.56 1.04 2.673 1.089 ;
      RECT 1.819 0.687 1.909 1.149 ;
      RECT 2.598 0.998 2.719 1.051 ;
      RECT 2.644 0.96 2.673 1.089 ;
      RECT 2.673 0.63 2.763 1.006 ;
      RECT 1.671 0.687 1.909 0.777 ;
      RECT 1.671 0.241 1.761 0.777 ;
      RECT 1.318 0.241 1.761 0.331 ;
      RECT 2.392 0.865 2.532 0.955 ;
      RECT 2.392 0.28 2.482 0.955 ;
      RECT 2.235 0.598 2.482 0.738 ;
      RECT 2.392 0.28 2.532 0.37 ;
      RECT 1.491 0.875 1.631 0.965 ;
      RECT 0.541 0.84 0.796 0.93 ;
      RECT 0.706 0.294 0.796 0.93 ;
      RECT 1.491 0.444 1.581 0.965 ;
      RECT 0.706 0.444 1.581 0.534 ;
      RECT 0.541 0.294 0.796 0.384 ;
      RECT 0.07 1.029 1.076 1.119 ;
      RECT 0.07 1.029 1.122 1.096 ;
      RECT 1.038 1.01 1.168 1.05 ;
      RECT 0.07 0.287 0.16 1.119 ;
      RECT 1.076 0.968 1.168 1.05 ;
      RECT 1.122 0.922 1.214 1.004 ;
      RECT 1.168 0.876 1.251 0.963 ;
      RECT 1.168 0.876 1.297 0.921 ;
      RECT 1.251 0.666 1.341 0.876 ;
      RECT 1.214 0.834 1.341 0.876 ;
      RECT 0.526 0.579 0.616 0.745 ;
      RECT 0.506 0.501 0.526 0.629 ;
      RECT 0.46 0.468 0.506 0.596 ;
      RECT 0.46 0.534 0.572 0.596 ;
      RECT 0.422 0.534 0.572 0.554 ;
      RECT 0.07 0.445 0.46 0.535 ;
  END
END LATHX1H7R

MACRO LATHX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATHX2H7R 0 0 ;
  SIZE 3.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.4 1.48 ;
        RECT 2.696 1.185 2.836 1.48 ;
        RECT 1.871 1.24 2.011 1.48 ;
        RECT 0.806 1.209 0.946 1.48 ;
        RECT 0.311 1.225 0.451 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.4 0.08 ;
        RECT 2.595 -0.08 2.685 0.335 ;
        RECT 1.851 -0.08 1.941 0.33 ;
        RECT 0.806 -0.08 0.946 0.204 ;
        RECT 0.295 -0.08 0.435 0.352 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.625 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.625 0.35 0.895 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END G
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.04 0.36 3.145 1.145 ;
        RECT 2.82 0.36 3.145 0.45 ;
      LAYER MET2 ;
        RECT 3.05 0.23 3.15 0.76 ;
      LAYER VIA1 ;
        RECT 3.055 0.455 3.145 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.055 0.83 2.341 0.92 ;
        RECT 2.055 0.36 2.216 0.45 ;
        RECT 2.055 0.36 2.145 0.92 ;
      LAYER MET2 ;
        RECT 2.05 0.23 2.15 0.76 ;
      LAYER VIA1 ;
        RECT 2.055 0.455 2.145 0.545 ;
    END
  END QN
  OBS
    LAYER MET1 ;
      RECT 1.301 1.059 2.602 1.149 ;
      RECT 2.564 1.04 2.682 1.092 ;
      RECT 2.602 1.004 2.636 1.132 ;
      RECT 1.819 0.687 1.909 1.149 ;
      RECT 2.636 0.62 2.726 1.047 ;
      RECT 1.671 0.687 1.909 0.777 ;
      RECT 2.636 0.62 2.926 0.76 ;
      RECT 1.671 0.241 1.761 0.777 ;
      RECT 1.318 0.241 1.761 0.331 ;
      RECT 2.456 0.598 2.546 0.945 ;
      RECT 2.235 0.598 2.546 0.738 ;
      RECT 2.345 0.255 2.435 0.738 ;
      RECT 1.481 0.879 1.621 0.969 ;
      RECT 0.541 0.84 0.796 0.93 ;
      RECT 0.706 0.294 0.796 0.93 ;
      RECT 1.481 0.465 1.571 0.969 ;
      RECT 1.222 0.465 1.571 0.555 ;
      RECT 1.181 0.406 1.222 0.535 ;
      RECT 1.135 0.363 1.181 0.491 ;
      RECT 1.135 0.446 1.26 0.491 ;
      RECT 1.089 0.317 1.135 0.445 ;
      RECT 1.051 0.363 1.181 0.403 ;
      RECT 0.541 0.294 1.089 0.384 ;
      RECT 0.07 1.029 1.076 1.119 ;
      RECT 0.07 1.029 1.122 1.096 ;
      RECT 1.038 1.01 1.168 1.05 ;
      RECT 0.07 0.287 0.16 1.119 ;
      RECT 1.076 0.968 1.168 1.05 ;
      RECT 1.214 0.84 1.24 0.968 ;
      RECT 1.122 0.922 1.24 0.968 ;
      RECT 1.168 0.876 1.214 1.004 ;
      RECT 1.24 0.666 1.286 0.932 ;
      RECT 1.24 0.666 1.33 0.887 ;
      RECT 0.526 0.569 0.616 0.745 ;
      RECT 0.516 0.496 0.526 0.624 ;
      RECT 0.47 0.468 0.516 0.596 ;
      RECT 0.47 0.524 0.572 0.596 ;
      RECT 0.432 0.524 0.572 0.554 ;
      RECT 0.07 0.445 0.47 0.535 ;
  END
END LATHX2H7R

MACRO LATHX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATHX3H7R 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.8 1.48 ;
        RECT 3.633 0.955 3.723 1.48 ;
        RECT 3.093 1.225 3.243 1.48 ;
        RECT 2.63 1.2 2.72 1.48 ;
        RECT 2.037 1.225 2.177 1.48 ;
        RECT 0.806 1.209 0.946 1.48 ;
        RECT 0.311 1.225 0.451 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.8 0.08 ;
        RECT 3.602 -0.08 3.692 0.345 ;
        RECT 3.102 -0.08 3.192 0.33 ;
        RECT 2.606 -0.08 2.696 0.35 ;
        RECT 2.045 -0.08 2.135 0.33 ;
        RECT 0.806 -0.08 0.946 0.204 ;
        RECT 0.295 -0.08 0.435 0.352 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.625 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.625 0.35 0.895 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END G
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.383 0.655 3.575 0.745 ;
        RECT 3.383 0.305 3.473 0.945 ;
        RECT 3.327 0.305 3.473 0.395 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.225 0.255 2.471 0.345 ;
        RECT 2.321 0.828 2.461 0.985 ;
        RECT 2.225 0.828 2.461 0.918 ;
        RECT 2.225 0.255 2.315 0.918 ;
      LAYER MET2 ;
        RECT 2.25 0.18 2.35 0.56 ;
      LAYER VIA1 ;
        RECT 2.255 0.255 2.345 0.345 ;
    END
  END QN
  OBS
    LAYER MET1 ;
      RECT 1.321 1.02 1.411 1.174 ;
      RECT 2.245 1.075 2.537 1.165 ;
      RECT 2.228 1.075 2.554 1.157 ;
      RECT 2.19 1.075 2.592 1.129 ;
      RECT 3.057 0.62 3.147 1.11 ;
      RECT 2.499 1.056 3.147 1.11 ;
      RECT 2.554 1.02 3.147 1.11 ;
      RECT 1.321 1.056 2.283 1.11 ;
      RECT 2.537 1.028 3.147 1.11 ;
      RECT 1.321 1.028 2.245 1.11 ;
      RECT 1.321 1.02 2.228 1.11 ;
      RECT 1.99 0.638 2.08 1.11 ;
      RECT 1.983 0.566 1.99 0.695 ;
      RECT 1.937 0.54 1.983 0.668 ;
      RECT 1.937 0.593 2.036 0.668 ;
      RECT 1.891 0.494 1.937 0.622 ;
      RECT 1.845 0.448 1.891 0.576 ;
      RECT 1.799 0.402 1.845 0.53 ;
      RECT 1.753 0.356 1.799 0.484 ;
      RECT 1.707 0.31 1.753 0.438 ;
      RECT 1.661 0.264 1.707 0.392 ;
      RECT 1.623 0.31 1.753 0.35 ;
      RECT 1.318 0.241 1.661 0.331 ;
      RECT 2.827 0.83 2.967 0.92 ;
      RECT 2.827 0.28 2.917 0.92 ;
      RECT 2.41 0.623 2.917 0.713 ;
      RECT 2.827 0.28 2.967 0.37 ;
      RECT 0.541 0.849 0.796 0.939 ;
      RECT 0.706 0.294 0.796 0.939 ;
      RECT 1.687 0.683 1.777 0.9 ;
      RECT 1.644 0.593 1.687 0.722 ;
      RECT 1.644 0.638 1.733 0.722 ;
      RECT 1.598 0.549 1.644 0.677 ;
      RECT 1.552 0.503 1.598 0.631 ;
      RECT 1.247 0.48 1.337 0.62 ;
      RECT 1.514 0.549 1.644 0.589 ;
      RECT 1.227 0.48 1.552 0.57 ;
      RECT 1.181 0.409 1.227 0.537 ;
      RECT 1.135 0.363 1.181 0.491 ;
      RECT 1.135 0.466 1.275 0.491 ;
      RECT 1.135 0.442 1.247 0.491 ;
      RECT 1.089 0.317 1.135 0.445 ;
      RECT 1.051 0.363 1.181 0.403 ;
      RECT 0.541 0.294 1.089 0.384 ;
      RECT 0.07 1.029 1.076 1.119 ;
      RECT 0.07 1.029 1.122 1.096 ;
      RECT 1.038 1.01 1.168 1.05 ;
      RECT 0.07 0.287 0.16 1.119 ;
      RECT 1.076 0.968 1.168 1.05 ;
      RECT 1.122 0.922 1.214 1.004 ;
      RECT 1.122 0.922 1.26 0.958 ;
      RECT 1.168 0.876 1.277 0.927 ;
      RECT 1.168 0.876 1.315 0.899 ;
      RECT 1.457 0.74 1.547 0.88 ;
      RECT 1.214 0.83 1.547 0.88 ;
      RECT 1.277 0.79 1.547 0.88 ;
      RECT 1.26 0.798 1.547 0.88 ;
      RECT 0.526 0.574 0.616 0.745 ;
      RECT 0.511 0.498 0.526 0.627 ;
      RECT 0.465 0.468 0.511 0.596 ;
      RECT 0.465 0.529 0.572 0.596 ;
      RECT 0.427 0.529 0.572 0.554 ;
      RECT 0.07 0.445 0.465 0.535 ;
  END
END LATHX3H7R

MACRO LATHX4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATHX4H7R 0 0 ;
  SIZE 4.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.4 1.48 ;
        RECT 3.933 1.035 4.073 1.48 ;
        RECT 3.403 1.225 3.543 1.48 ;
        RECT 2.612 1.24 2.752 1.48 ;
        RECT 2.037 1.225 2.177 1.48 ;
        RECT 0.821 1.224 0.961 1.48 ;
        RECT 0.311 1.225 0.451 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.4 0.08 ;
        RECT 3.572 -0.08 3.712 0.34 ;
        RECT 3.097 -0.08 3.187 0.35 ;
        RECT 2.606 -0.08 2.696 0.35 ;
        RECT 2.045 -0.08 2.135 0.33 ;
        RECT 0.806 -0.08 0.946 0.204 ;
        RECT 0.295 -0.08 0.435 0.352 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.625 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.625 0.35 0.895 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END G
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.668 0.855 4.338 0.945 ;
        RECT 4.248 0.465 4.338 0.945 ;
        RECT 3.347 0.465 4.338 0.555 ;
        RECT 3.347 0.37 3.437 0.555 ;
      LAYER MET2 ;
        RECT 3.85 0.63 3.95 1.16 ;
      LAYER VIA1 ;
        RECT 3.855 0.855 3.945 0.945 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.892 0.855 3.032 0.985 ;
        RECT 2.321 0.855 3.032 0.945 ;
        RECT 2.321 0.375 2.471 0.465 ;
        RECT 2.321 0.855 2.461 0.985 ;
        RECT 2.321 0.375 2.411 0.985 ;
      LAYER MET2 ;
        RECT 2.45 0.625 2.55 1.16 ;
      LAYER VIA1 ;
        RECT 2.455 0.855 2.545 0.945 ;
    END
  END QN
  OBS
    LAYER MET1 ;
      RECT 2.514 1.06 2.517 1.185 ;
      RECT 2.303 1.095 2.479 1.185 ;
      RECT 2.843 1.075 3.271 1.165 ;
      RECT 2.805 1.06 2.828 1.165 ;
      RECT 2.552 1.06 2.79 1.15 ;
      RECT 2.08 1.045 2.215 1.135 ;
      RECT 1.562 1.045 1.99 1.135 ;
      RECT 3.432 0.645 4.082 0.735 ;
      RECT 1.318 0.241 1.623 0.331 ;
      RECT 3.388 0.645 3.432 1.064 ;
      RECT 3.342 0.645 3.388 1.109 ;
      RECT 3.309 1.02 3.342 1.149 ;
      RECT 3.271 1.056 3.309 1.165 ;
      RECT 2.828 1.067 2.843 1.165 ;
      RECT 2.79 1.06 2.805 1.158 ;
      RECT 2.517 1.06 2.552 1.168 ;
      RECT 2.479 1.077 2.514 1.185 ;
      RECT 2.265 1.076 2.303 1.185 ;
      RECT 2.253 1.051 2.265 1.179 ;
      RECT 2.215 1.045 2.253 1.154 ;
      RECT 2.036 0.638 2.08 1.135 ;
      RECT 1.99 0.593 2.036 1.135 ;
      RECT 1.983 0.566 1.99 0.695 ;
      RECT 1.937 0.54 1.983 0.668 ;
      RECT 1.891 0.494 1.937 0.622 ;
      RECT 1.845 0.448 1.891 0.576 ;
      RECT 1.799 0.402 1.845 0.53 ;
      RECT 1.753 0.356 1.799 0.484 ;
      RECT 1.707 0.31 1.753 0.438 ;
      RECT 1.661 0.264 1.707 0.392 ;
      RECT 1.623 0.241 1.661 0.35 ;
      RECT 3.162 0.623 3.252 0.965 ;
      RECT 2.512 0.623 3.252 0.713 ;
      RECT 2.847 0.255 2.937 0.713 ;
      RECT 0.541 0.849 0.796 0.939 ;
      RECT 0.706 0.294 0.796 0.939 ;
      RECT 1.687 0.683 1.777 0.9 ;
      RECT 1.644 0.593 1.687 0.722 ;
      RECT 1.644 0.638 1.733 0.722 ;
      RECT 1.598 0.549 1.644 0.677 ;
      RECT 1.552 0.503 1.598 0.631 ;
      RECT 1.247 0.48 1.337 0.62 ;
      RECT 1.514 0.549 1.644 0.589 ;
      RECT 1.227 0.48 1.552 0.57 ;
      RECT 1.181 0.409 1.227 0.537 ;
      RECT 1.135 0.363 1.181 0.491 ;
      RECT 1.135 0.466 1.275 0.491 ;
      RECT 1.135 0.442 1.247 0.491 ;
      RECT 1.089 0.317 1.135 0.445 ;
      RECT 1.051 0.363 1.181 0.403 ;
      RECT 0.541 0.294 1.089 0.384 ;
      RECT 0.07 1.029 1.076 1.119 ;
      RECT 0.07 1.029 1.122 1.096 ;
      RECT 1.038 1.01 1.168 1.05 ;
      RECT 0.07 0.287 0.16 1.119 ;
      RECT 1.076 0.968 1.168 1.05 ;
      RECT 1.122 0.922 1.214 1.004 ;
      RECT 1.122 0.922 1.26 0.958 ;
      RECT 1.168 0.876 1.277 0.927 ;
      RECT 1.168 0.876 1.315 0.899 ;
      RECT 1.457 0.74 1.547 0.88 ;
      RECT 1.214 0.83 1.547 0.88 ;
      RECT 1.277 0.79 1.547 0.88 ;
      RECT 1.26 0.798 1.547 0.88 ;
      RECT 0.526 0.574 0.616 0.745 ;
      RECT 0.511 0.498 0.526 0.627 ;
      RECT 0.465 0.468 0.511 0.596 ;
      RECT 0.465 0.529 0.572 0.596 ;
      RECT 0.427 0.529 0.572 0.554 ;
      RECT 0.07 0.445 0.465 0.535 ;
  END
END LATHX4H7R

MACRO LATLRX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATLRX0P5H7R 0 0 ;
  SIZE 4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4 1.48 ;
        RECT 3.52 1.055 3.61 1.48 ;
        RECT 2.8 1.07 2.89 1.48 ;
        RECT 2.32 1.035 2.41 1.48 ;
        RECT 1.555 1.24 1.695 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4 0.08 ;
        RECT 3.51 -0.08 3.6 0.33 ;
        RECT 3.015 -0.08 3.105 0.33 ;
        RECT 1.76 -0.08 1.9 0.175 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.44 0.565 1.56 0.79 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.715 0.375 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END GN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.16 0.405 3.355 0.495 ;
        RECT 3.255 0.225 3.355 0.495 ;
        RECT 3.16 0.405 3.25 1.05 ;
      LAYER MET2 ;
        RECT 3.25 0.18 3.35 0.56 ;
      LAYER VIA1 ;
        RECT 3.255 0.255 3.345 0.345 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.77 0.425 3.945 0.575 ;
        RECT 3.77 0.255 3.86 1.065 ;
      LAYER MET2 ;
        RECT 3.85 0.23 3.95 0.76 ;
      LAYER VIA1 ;
        RECT 3.855 0.455 3.945 0.545 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.75 0.455 1.975 0.575 ;
      LAYER MET2 ;
        RECT 1.85 0.225 1.95 0.76 ;
      LAYER VIA1 ;
        RECT 1.855 0.455 1.945 0.545 ;
    END
  END RN
  OBS
    LAYER MET1 ;
      RECT 2.98 1.14 3.43 1.23 ;
      RECT 3.34 0.765 3.43 1.23 ;
      RECT 2.98 0.42 3.07 1.23 ;
      RECT 2.525 0.855 2.665 1.04 ;
      RECT 2.32 0.855 3.07 0.945 ;
      RECT 3.34 0.765 3.68 0.855 ;
      RECT 3.59 0.715 3.68 0.855 ;
      RECT 2.32 0.805 2.41 0.945 ;
      RECT 2.765 0.42 3.07 0.51 ;
      RECT 2.765 0.255 2.855 0.51 ;
      RECT 0.86 1.13 1.29 1.22 ;
      RECT 0.86 1.13 1.321 1.205 ;
      RECT 0.86 1.13 1.36 1.17 ;
      RECT 2.14 0.625 2.23 1.15 ;
      RECT 1.251 1.11 2.23 1.15 ;
      RECT 1.321 1.06 2.23 1.15 ;
      RECT 0.86 0.35 0.95 1.22 ;
      RECT 1.29 1.075 2.23 1.15 ;
      RECT 0.825 0.948 0.95 1.088 ;
      RECT 2.14 0.625 2.845 0.715 ;
      RECT 2.585 0.25 2.675 0.715 ;
      RECT 0.79 0.35 0.95 0.44 ;
      RECT 2.51 0.25 2.675 0.34 ;
      RECT 0.545 0.95 0.7 1.04 ;
      RECT 0.61 0.17 0.7 1.04 ;
      RECT 0.61 0.688 0.77 0.828 ;
      RECT 2.139 0.435 2.485 0.525 ;
      RECT 2.139 0.265 2.229 0.525 ;
      RECT 1.497 0.265 2.229 0.355 ;
      RECT 1.487 0.221 1.497 0.35 ;
      RECT 0.57 0.17 0.7 0.348 ;
      RECT 1.441 0.193 1.487 0.322 ;
      RECT 1.402 0.245 1.536 0.28 ;
      RECT 0.57 0.17 1.441 0.26 ;
      RECT 1.255 0.88 2.05 0.97 ;
      RECT 1.96 0.775 2.05 0.97 ;
      RECT 1.255 0.555 1.345 0.97 ;
      RECT 1.22 0.555 1.345 0.695 ;
      RECT 1.04 0.9 1.165 1.04 ;
      RECT 1.04 0.35 1.13 1.04 ;
      RECT 1.04 0.35 1.24 0.44 ;
      RECT 0.045 1.01 0.16 1.15 ;
      RECT 0.045 0.28 0.135 1.15 ;
      RECT 0.43 0.465 0.52 0.605 ;
      RECT 0.045 0.465 0.52 0.555 ;
      RECT 0.045 0.28 0.185 0.37 ;
  END
END LATLRX0P5H7R

MACRO LATLRX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATLRX1H7R 0 0 ;
  SIZE 4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4 1.48 ;
        RECT 3.52 1.055 3.61 1.48 ;
        RECT 2.8 1.07 2.89 1.48 ;
        RECT 2.32 1.035 2.41 1.48 ;
        RECT 1.555 1.24 1.695 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4 0.08 ;
        RECT 3.51 -0.08 3.6 0.33 ;
        RECT 3.015 -0.08 3.105 0.33 ;
        RECT 1.76 -0.08 1.9 0.175 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.44 0.565 1.56 0.79 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.715 0.375 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END GN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.16 0.485 3.355 0.575 ;
        RECT 3.255 0.295 3.355 0.575 ;
        RECT 3.16 0.485 3.25 1.005 ;
      LAYER MET2 ;
        RECT 3.25 0.23 3.35 0.76 ;
      LAYER VIA1 ;
        RECT 3.255 0.455 3.345 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.77 0.425 3.945 0.575 ;
        RECT 3.77 0.295 3.86 1.005 ;
      LAYER MET2 ;
        RECT 3.85 0.23 3.95 0.76 ;
      LAYER VIA1 ;
        RECT 3.855 0.455 3.945 0.545 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.75 0.455 1.975 0.575 ;
      LAYER MET2 ;
        RECT 1.85 0.225 1.95 0.76 ;
      LAYER VIA1 ;
        RECT 1.855 0.455 1.945 0.545 ;
    END
  END RN
  OBS
    LAYER MET1 ;
      RECT 2.98 1.095 3.43 1.185 ;
      RECT 3.34 0.705 3.43 1.185 ;
      RECT 2.98 0.42 3.07 1.185 ;
      RECT 2.525 0.855 2.665 1.04 ;
      RECT 2.32 0.855 3.07 0.945 ;
      RECT 2.32 0.805 2.41 0.945 ;
      RECT 3.34 0.705 3.68 0.795 ;
      RECT 3.59 0.655 3.68 0.795 ;
      RECT 2.765 0.42 3.07 0.51 ;
      RECT 2.765 0.255 2.855 0.51 ;
      RECT 0.86 1.14 1.28 1.23 ;
      RECT 0.86 1.14 1.321 1.21 ;
      RECT 0.86 1.14 1.36 1.17 ;
      RECT 2.14 0.625 2.23 1.15 ;
      RECT 1.241 1.12 2.23 1.15 ;
      RECT 1.321 1.06 2.23 1.15 ;
      RECT 0.86 0.35 0.95 1.23 ;
      RECT 1.28 1.08 2.23 1.15 ;
      RECT 0.825 0.948 0.95 1.088 ;
      RECT 2.14 0.625 2.845 0.715 ;
      RECT 2.585 0.25 2.675 0.715 ;
      RECT 0.79 0.35 0.95 0.44 ;
      RECT 2.51 0.25 2.675 0.34 ;
      RECT 0.545 0.95 0.7 1.04 ;
      RECT 0.61 0.17 0.7 1.04 ;
      RECT 0.61 0.688 0.77 0.828 ;
      RECT 2.139 0.435 2.485 0.525 ;
      RECT 2.139 0.265 2.229 0.525 ;
      RECT 1.497 0.265 2.229 0.355 ;
      RECT 1.487 0.221 1.497 0.35 ;
      RECT 0.57 0.17 0.7 0.348 ;
      RECT 1.441 0.193 1.487 0.322 ;
      RECT 1.402 0.245 1.536 0.28 ;
      RECT 0.57 0.17 1.441 0.26 ;
      RECT 1.255 0.88 2.05 0.97 ;
      RECT 1.96 0.775 2.05 0.97 ;
      RECT 1.255 0.555 1.345 0.97 ;
      RECT 1.22 0.555 1.345 0.695 ;
      RECT 1.04 0.91 1.165 1.05 ;
      RECT 1.04 0.35 1.13 1.05 ;
      RECT 1.04 0.35 1.24 0.44 ;
      RECT 0.045 1.01 0.16 1.15 ;
      RECT 0.045 0.28 0.135 1.15 ;
      RECT 0.43 0.465 0.52 0.605 ;
      RECT 0.045 0.465 0.52 0.555 ;
      RECT 0.045 0.28 0.185 0.37 ;
  END
END LATLRX1H7R

MACRO LATLRX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATLRX2H7R 0 0 ;
  SIZE 4.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.2 1.48 ;
        RECT 4.02 1.052 4.11 1.48 ;
        RECT 3.52 1.07 3.61 1.48 ;
        RECT 2.8 1.07 2.89 1.48 ;
        RECT 2.32 1.035 2.41 1.48 ;
        RECT 1.555 1.24 1.695 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.2 0.08 ;
        RECT 4.02 -0.08 4.11 0.341 ;
        RECT 3.51 -0.08 3.6 0.33 ;
        RECT 3.015 -0.08 3.105 0.33 ;
        RECT 1.76 -0.08 1.9 0.175 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.44 0.565 1.56 0.79 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.715 0.375 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END GN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.16 0.485 3.355 0.575 ;
        RECT 3.255 0.335 3.355 0.575 ;
        RECT 3.16 0.485 3.25 1.05 ;
      LAYER MET2 ;
        RECT 3.25 0.23 3.35 0.76 ;
      LAYER VIA1 ;
        RECT 3.255 0.455 3.345 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.77 0.425 3.945 0.575 ;
        RECT 3.77 0.21 3.86 1.13 ;
      LAYER MET2 ;
        RECT 3.85 0.23 3.95 0.76 ;
      LAYER VIA1 ;
        RECT 3.855 0.455 3.945 0.545 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.75 0.455 1.975 0.575 ;
      LAYER MET2 ;
        RECT 1.85 0.225 1.95 0.76 ;
      LAYER VIA1 ;
        RECT 1.855 0.455 1.945 0.545 ;
    END
  END RN
  OBS
    LAYER MET1 ;
      RECT 2.98 1.14 3.43 1.23 ;
      RECT 3.34 0.795 3.43 1.23 ;
      RECT 2.98 0.42 3.07 1.23 ;
      RECT 2.525 0.855 2.665 1.04 ;
      RECT 2.32 0.855 3.07 0.945 ;
      RECT 3.34 0.795 3.68 0.935 ;
      RECT 2.32 0.805 2.41 0.945 ;
      RECT 2.765 0.42 3.07 0.51 ;
      RECT 2.765 0.255 2.855 0.51 ;
      RECT 0.86 1.14 1.28 1.23 ;
      RECT 0.86 1.14 1.321 1.21 ;
      RECT 0.86 1.14 1.36 1.17 ;
      RECT 2.14 0.625 2.23 1.15 ;
      RECT 1.241 1.12 2.23 1.15 ;
      RECT 1.321 1.06 2.23 1.15 ;
      RECT 0.86 0.35 0.95 1.23 ;
      RECT 1.28 1.08 2.23 1.15 ;
      RECT 0.825 0.948 0.95 1.088 ;
      RECT 2.14 0.625 2.845 0.715 ;
      RECT 2.585 0.25 2.675 0.715 ;
      RECT 0.79 0.35 0.95 0.44 ;
      RECT 2.51 0.25 2.675 0.34 ;
      RECT 0.545 0.95 0.7 1.04 ;
      RECT 0.61 0.17 0.7 1.04 ;
      RECT 0.61 0.688 0.77 0.828 ;
      RECT 2.139 0.435 2.485 0.525 ;
      RECT 2.139 0.265 2.229 0.525 ;
      RECT 1.497 0.265 2.229 0.355 ;
      RECT 1.487 0.221 1.497 0.35 ;
      RECT 0.57 0.17 0.7 0.348 ;
      RECT 1.441 0.193 1.487 0.322 ;
      RECT 1.402 0.245 1.536 0.28 ;
      RECT 0.57 0.17 1.441 0.26 ;
      RECT 1.255 0.88 2.05 0.97 ;
      RECT 1.96 0.775 2.05 0.97 ;
      RECT 1.255 0.555 1.345 0.97 ;
      RECT 1.22 0.555 1.345 0.695 ;
      RECT 1.04 0.91 1.165 1.05 ;
      RECT 1.04 0.35 1.13 1.05 ;
      RECT 1.04 0.35 1.24 0.44 ;
      RECT 0.045 1.01 0.16 1.15 ;
      RECT 0.045 0.28 0.135 1.15 ;
      RECT 0.43 0.465 0.52 0.605 ;
      RECT 0.045 0.465 0.52 0.555 ;
      RECT 0.045 0.28 0.185 0.37 ;
  END
END LATLRX2H7R

MACRO LATLSRX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATLSRX0P5H7R 0 0 ;
  SIZE 6.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.8 1.48 ;
        RECT 6.245 1.07 6.335 1.48 ;
        RECT 5.125 1.24 5.265 1.48 ;
        RECT 4.244 1.095 4.384 1.48 ;
        RECT 0.325 1.095 0.465 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.8 0.08 ;
        RECT 6.195 -0.08 6.335 0.16 ;
        RECT 5.125 -0.08 5.265 0.16 ;
        RECT 4.119 -0.08 4.209 0.33 ;
        RECT 0.375 -0.08 0.465 0.33 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.843 0.735 3.145 0.825 ;
        RECT 3.055 0.625 3.145 0.825 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.655 0.385 0.825 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END GN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.865 0.36 6.005 0.45 ;
        RECT 5.825 0.855 5.975 0.965 ;
        RECT 5.865 0.36 5.955 0.965 ;
      LAYER MET2 ;
        RECT 5.85 0.63 5.95 1.16 ;
      LAYER VIA1 ;
        RECT 5.855 0.855 5.945 0.945 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.455 0.875 5.595 0.965 ;
        RECT 5.455 0.36 5.595 0.45 ;
        RECT 5.455 0.36 5.545 0.965 ;
      LAYER MET2 ;
        RECT 5.45 0.225 5.55 0.76 ;
      LAYER VIA1 ;
        RECT 5.455 0.455 5.545 0.545 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.03 0.42 4.15 0.645 ;
      LAYER MET2 ;
        RECT 4.05 0.23 4.15 0.76 ;
      LAYER VIA1 ;
        RECT 4.055 0.455 4.145 0.545 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.975 0.625 5.155 0.775 ;
      LAYER MET2 ;
        RECT 5.05 0.43 5.15 0.96 ;
      LAYER VIA1 ;
        RECT 5.055 0.655 5.145 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 6.55 0.255 6.64 1.065 ;
      RECT 3.85 0.735 4.389 0.825 ;
      RECT 4.299 0.17 4.389 0.825 ;
      RECT 3.85 0.45 3.94 0.825 ;
      RECT 5.685 0.17 5.775 0.666 ;
      RECT 3.499 0.45 3.94 0.54 ;
      RECT 6.119 0.255 6.64 0.345 ;
      RECT 5.022 0.25 5.341 0.34 ;
      RECT 6.073 0.193 6.119 0.321 ;
      RECT 4.98 0.25 5.383 0.319 ;
      RECT 6.035 0.255 6.64 0.279 ;
      RECT 4.942 0.25 5.421 0.279 ;
      RECT 5.383 0.17 6.073 0.26 ;
      RECT 6.119 0.236 6.158 0.345 ;
      RECT 5.341 0.191 5.383 0.319 ;
      RECT 4.299 0.231 5.06 0.26 ;
      RECT 5.303 0.231 6.12 0.26 ;
      RECT 6.119 0.216 6.12 0.345 ;
      RECT 4.299 0.191 5.022 0.26 ;
      RECT 4.299 0.17 4.98 0.26 ;
      RECT 4.48 1.06 6.155 1.15 ;
      RECT 6.065 0.572 6.155 1.15 ;
      RECT 4.48 0.35 4.57 1.15 ;
      RECT 3.67 0.915 3.81 1.05 ;
      RECT 3.67 0.915 4.57 1.005 ;
      RECT 1.13 0.865 1.249 1.005 ;
      RECT 1.159 0.17 1.249 1.005 ;
      RECT 3.67 0.645 3.76 1.05 ;
      RECT 3.438 0.645 3.76 0.735 ;
      RECT 3.426 0.601 3.438 0.729 ;
      RECT 3.38 0.572 3.426 0.7 ;
      RECT 6.065 0.572 6.405 0.662 ;
      RECT 3.334 0.526 3.38 0.654 ;
      RECT 3.334 0.626 3.476 0.654 ;
      RECT 3.288 0.48 3.334 0.608 ;
      RECT 3.242 0.434 3.288 0.562 ;
      RECT 3.196 0.388 3.242 0.516 ;
      RECT 3.158 0.434 3.288 0.474 ;
      RECT 2.149 0.365 3.196 0.455 ;
      RECT 4.48 0.35 4.62 0.44 ;
      RECT 1.629 0.17 1.769 0.367 ;
      RECT 2.149 0.17 2.239 0.455 ;
      RECT 1.159 0.17 2.239 0.26 ;
      RECT 4.71 0.876 4.85 0.97 ;
      RECT 4.71 0.35 4.8 0.97 ;
      RECT 4.71 0.35 4.88 0.44 ;
      RECT 1.9 1.14 4.134 1.23 ;
      RECT 3.994 1.095 4.134 1.23 ;
      RECT 3.08 1.095 3.22 1.23 ;
      RECT 3.416 0.215 3.984 0.305 ;
      RECT 2.329 0.185 3.505 0.275 ;
      RECT 2.475 0.915 3.58 1.005 ;
      RECT 3.44 0.895 3.58 1.005 ;
      RECT 2.475 0.78 2.565 1.005 ;
      RECT 1.739 0.78 2.565 0.87 ;
      RECT 1.739 0.65 1.879 0.87 ;
      RECT 1.38 1.06 1.8 1.15 ;
      RECT 1.71 0.96 1.8 1.15 ;
      RECT 1.38 0.829 1.47 1.15 ;
      RECT 1.71 0.96 2.385 1.05 ;
      RECT 1.339 0.37 1.429 0.868 ;
      RECT 1.969 0.545 2.779 0.635 ;
      RECT 1.339 0.457 2.059 0.547 ;
      RECT 1.969 0.37 2.059 0.635 ;
      RECT 0.555 1.14 1.04 1.23 ;
      RECT 0.95 0.475 1.04 1.23 ;
      RECT 0.555 0.915 0.645 1.23 ;
      RECT 0.045 0.915 0.19 1.065 ;
      RECT 0.045 0.915 0.645 1.005 ;
      RECT 0.045 0.28 0.135 1.065 ;
      RECT 0.47 0.471 0.56 0.62 ;
      RECT 0.95 0.475 1.069 0.615 ;
      RECT 0.045 0.471 0.56 0.561 ;
      RECT 0.045 0.28 0.215 0.37 ;
      RECT 0.735 0.28 0.825 1.05 ;
      RECT 0.6 0.28 0.825 0.37 ;
  END
END LATLSRX0P5H7R

MACRO LATLSRX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATLSRX1H7R 0 0 ;
  SIZE 6.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.8 1.48 ;
        RECT 6.245 1.07 6.335 1.48 ;
        RECT 5.125 1.24 5.265 1.48 ;
        RECT 4.244 1.095 4.384 1.48 ;
        RECT 0.325 1.095 0.465 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.8 0.08 ;
        RECT 6.195 -0.08 6.335 0.16 ;
        RECT 5.125 -0.08 5.265 0.16 ;
        RECT 4.119 -0.08 4.209 0.33 ;
        RECT 0.375 -0.08 0.465 0.33 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.843 0.735 3.145 0.825 ;
        RECT 3.055 0.625 3.145 0.825 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.655 0.385 0.825 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END GN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.865 0.36 6.005 0.45 ;
        RECT 5.825 0.855 5.975 0.965 ;
        RECT 5.865 0.36 5.955 0.965 ;
      LAYER MET2 ;
        RECT 5.85 0.63 5.95 1.16 ;
      LAYER VIA1 ;
        RECT 5.855 0.855 5.945 0.945 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.455 0.875 5.595 0.965 ;
        RECT 5.455 0.36 5.595 0.45 ;
        RECT 5.455 0.36 5.545 0.965 ;
      LAYER MET2 ;
        RECT 5.45 0.225 5.55 0.76 ;
      LAYER VIA1 ;
        RECT 5.455 0.455 5.545 0.545 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.03 0.42 4.15 0.645 ;
      LAYER MET2 ;
        RECT 4.05 0.23 4.15 0.76 ;
      LAYER VIA1 ;
        RECT 4.055 0.455 4.145 0.545 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.975 0.625 5.155 0.775 ;
      LAYER MET2 ;
        RECT 5.05 0.43 5.15 0.96 ;
      LAYER VIA1 ;
        RECT 5.055 0.655 5.145 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 6.55 0.255 6.64 1.065 ;
      RECT 3.85 0.735 4.389 0.825 ;
      RECT 4.299 0.17 4.389 0.825 ;
      RECT 3.85 0.45 3.94 0.825 ;
      RECT 5.685 0.17 5.775 0.666 ;
      RECT 3.499 0.45 3.94 0.54 ;
      RECT 6.119 0.255 6.64 0.345 ;
      RECT 5.022 0.25 5.341 0.34 ;
      RECT 6.073 0.193 6.119 0.321 ;
      RECT 4.98 0.25 5.383 0.319 ;
      RECT 6.035 0.255 6.64 0.279 ;
      RECT 4.942 0.25 5.421 0.279 ;
      RECT 5.383 0.17 6.073 0.26 ;
      RECT 6.119 0.236 6.158 0.345 ;
      RECT 5.341 0.191 5.383 0.319 ;
      RECT 4.299 0.231 5.06 0.26 ;
      RECT 5.303 0.231 6.12 0.26 ;
      RECT 6.119 0.216 6.12 0.345 ;
      RECT 4.299 0.191 5.022 0.26 ;
      RECT 4.299 0.17 4.98 0.26 ;
      RECT 4.48 1.06 6.155 1.15 ;
      RECT 6.065 0.572 6.155 1.15 ;
      RECT 4.48 0.35 4.57 1.15 ;
      RECT 3.67 0.915 3.81 1.05 ;
      RECT 3.67 0.915 4.57 1.005 ;
      RECT 1.13 0.865 1.249 1.005 ;
      RECT 1.159 0.17 1.249 1.005 ;
      RECT 3.67 0.645 3.76 1.05 ;
      RECT 3.438 0.645 3.76 0.735 ;
      RECT 3.426 0.601 3.438 0.729 ;
      RECT 3.38 0.572 3.426 0.7 ;
      RECT 6.065 0.572 6.405 0.662 ;
      RECT 3.334 0.526 3.38 0.654 ;
      RECT 3.334 0.626 3.476 0.654 ;
      RECT 3.288 0.48 3.334 0.608 ;
      RECT 3.242 0.434 3.288 0.562 ;
      RECT 3.196 0.388 3.242 0.516 ;
      RECT 3.158 0.434 3.288 0.474 ;
      RECT 2.149 0.365 3.196 0.455 ;
      RECT 4.48 0.35 4.62 0.44 ;
      RECT 1.629 0.17 1.769 0.367 ;
      RECT 2.149 0.17 2.239 0.455 ;
      RECT 1.159 0.17 2.239 0.26 ;
      RECT 4.71 0.876 4.85 0.97 ;
      RECT 4.71 0.35 4.8 0.97 ;
      RECT 4.71 0.35 4.88 0.44 ;
      RECT 1.9 1.14 4.134 1.23 ;
      RECT 3.994 1.095 4.134 1.23 ;
      RECT 3.08 1.095 3.22 1.23 ;
      RECT 3.416 0.215 3.984 0.305 ;
      RECT 2.329 0.185 3.505 0.275 ;
      RECT 2.475 0.915 3.58 1.005 ;
      RECT 3.44 0.895 3.58 1.005 ;
      RECT 2.475 0.78 2.565 1.005 ;
      RECT 1.739 0.78 2.565 0.87 ;
      RECT 1.739 0.65 1.879 0.87 ;
      RECT 1.38 1.06 1.8 1.15 ;
      RECT 1.71 0.96 1.8 1.15 ;
      RECT 1.38 0.829 1.47 1.15 ;
      RECT 1.71 0.96 2.385 1.05 ;
      RECT 1.339 0.37 1.429 0.868 ;
      RECT 1.969 0.545 2.779 0.635 ;
      RECT 1.339 0.457 2.059 0.547 ;
      RECT 1.969 0.37 2.059 0.635 ;
      RECT 0.555 1.14 1.04 1.23 ;
      RECT 0.95 0.475 1.04 1.23 ;
      RECT 0.555 0.915 0.645 1.23 ;
      RECT 0.045 0.915 0.19 1.065 ;
      RECT 0.045 0.915 0.645 1.005 ;
      RECT 0.045 0.28 0.135 1.065 ;
      RECT 0.47 0.471 0.56 0.62 ;
      RECT 0.95 0.475 1.069 0.615 ;
      RECT 0.045 0.471 0.56 0.561 ;
      RECT 0.045 0.28 0.215 0.37 ;
      RECT 0.735 0.28 0.825 1.05 ;
      RECT 0.6 0.28 0.825 0.37 ;
  END
END LATLSRX1H7R

MACRO LATLSRX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATLSRX2H7R 0 0 ;
  SIZE 6.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.8 1.48 ;
        RECT 6.245 1.07 6.335 1.48 ;
        RECT 5.125 1.24 5.265 1.48 ;
        RECT 4.244 1.095 4.384 1.48 ;
        RECT 0.325 1.095 0.465 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.8 0.08 ;
        RECT 6.195 -0.08 6.335 0.16 ;
        RECT 5.125 -0.08 5.265 0.16 ;
        RECT 4.119 -0.08 4.209 0.33 ;
        RECT 0.375 -0.08 0.465 0.33 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.843 0.735 3.145 0.825 ;
        RECT 3.055 0.625 3.145 0.825 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.655 0.385 0.825 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END GN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.865 0.36 6.005 0.45 ;
        RECT 5.825 0.855 5.975 0.945 ;
        RECT 5.865 0.36 5.955 0.945 ;
      LAYER MET2 ;
        RECT 5.85 0.63 5.95 1.16 ;
      LAYER VIA1 ;
        RECT 5.855 0.855 5.945 0.945 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.455 0.83 5.595 0.92 ;
        RECT 5.455 0.36 5.595 0.45 ;
        RECT 5.455 0.36 5.545 0.92 ;
      LAYER MET2 ;
        RECT 5.45 0.225 5.55 0.76 ;
      LAYER VIA1 ;
        RECT 5.455 0.455 5.545 0.545 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.03 0.42 4.15 0.645 ;
      LAYER MET2 ;
        RECT 4.05 0.23 4.15 0.76 ;
      LAYER VIA1 ;
        RECT 4.055 0.455 4.145 0.545 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.975 0.625 5.155 0.775 ;
      LAYER MET2 ;
        RECT 5.05 0.43 5.15 0.96 ;
      LAYER VIA1 ;
        RECT 5.055 0.655 5.145 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 6.55 0.255 6.64 1.065 ;
      RECT 3.85 0.735 4.389 0.825 ;
      RECT 4.299 0.17 4.389 0.825 ;
      RECT 3.85 0.405 3.94 0.825 ;
      RECT 5.685 0.17 5.775 0.666 ;
      RECT 3.604 0.405 3.94 0.495 ;
      RECT 6.119 0.255 6.64 0.345 ;
      RECT 5.022 0.25 5.341 0.34 ;
      RECT 6.073 0.193 6.119 0.321 ;
      RECT 4.98 0.25 5.383 0.319 ;
      RECT 6.035 0.255 6.64 0.279 ;
      RECT 4.942 0.25 5.421 0.279 ;
      RECT 5.383 0.17 6.073 0.26 ;
      RECT 6.119 0.236 6.158 0.345 ;
      RECT 5.341 0.191 5.383 0.319 ;
      RECT 4.299 0.231 5.06 0.26 ;
      RECT 5.303 0.231 6.12 0.26 ;
      RECT 6.119 0.216 6.12 0.345 ;
      RECT 4.299 0.191 5.022 0.26 ;
      RECT 4.299 0.17 4.98 0.26 ;
      RECT 4.48 1.06 6.155 1.15 ;
      RECT 6.065 0.572 6.155 1.15 ;
      RECT 4.48 0.35 4.57 1.15 ;
      RECT 3.67 0.915 3.81 1.05 ;
      RECT 3.67 0.915 4.57 1.005 ;
      RECT 1.13 0.865 1.249 1.005 ;
      RECT 1.159 0.17 1.249 1.005 ;
      RECT 3.67 0.585 3.76 1.05 ;
      RECT 3.438 0.585 3.76 0.675 ;
      RECT 6.065 0.572 6.405 0.662 ;
      RECT 3.394 0.525 3.438 0.653 ;
      RECT 3.348 0.48 3.394 0.608 ;
      RECT 3.348 0.566 3.476 0.608 ;
      RECT 3.302 0.434 3.348 0.562 ;
      RECT 3.256 0.388 3.302 0.516 ;
      RECT 3.218 0.434 3.348 0.474 ;
      RECT 2.149 0.365 3.256 0.455 ;
      RECT 4.48 0.35 4.62 0.44 ;
      RECT 1.629 0.17 1.769 0.367 ;
      RECT 2.149 0.17 2.239 0.455 ;
      RECT 1.159 0.17 2.239 0.26 ;
      RECT 4.71 0.876 4.85 0.97 ;
      RECT 4.71 0.35 4.8 0.97 ;
      RECT 4.71 0.35 4.88 0.44 ;
      RECT 1.9 1.14 4.134 1.23 ;
      RECT 3.994 1.095 4.134 1.23 ;
      RECT 3.08 1.095 3.22 1.23 ;
      RECT 3.416 0.215 3.984 0.305 ;
      RECT 2.329 0.185 3.505 0.275 ;
      RECT 2.475 0.915 3.58 1.005 ;
      RECT 3.44 0.765 3.58 1.005 ;
      RECT 2.475 0.78 2.565 1.005 ;
      RECT 1.56 0.78 2.565 0.87 ;
      RECT 1.56 0.65 1.7 0.87 ;
      RECT 1.38 1.121 1.7 1.211 ;
      RECT 1.61 0.96 1.7 1.211 ;
      RECT 1.38 0.829 1.47 1.211 ;
      RECT 1.61 0.96 2.385 1.05 ;
      RECT 1.339 0.37 1.429 0.868 ;
      RECT 1.969 0.545 2.779 0.635 ;
      RECT 1.339 0.457 2.059 0.547 ;
      RECT 1.969 0.37 2.059 0.635 ;
      RECT 0.555 1.11 1.04 1.2 ;
      RECT 0.95 0.475 1.04 1.2 ;
      RECT 0.555 0.915 0.645 1.2 ;
      RECT 0.045 0.915 0.19 1.065 ;
      RECT 0.045 0.915 0.645 1.005 ;
      RECT 0.045 0.28 0.135 1.065 ;
      RECT 0.47 0.471 0.56 0.62 ;
      RECT 0.95 0.475 1.069 0.615 ;
      RECT 0.045 0.471 0.56 0.561 ;
      RECT 0.045 0.28 0.215 0.37 ;
      RECT 0.735 0.29 0.825 1.02 ;
      RECT 0.6 0.29 0.825 0.38 ;
  END
END LATLSRX2H7R

MACRO LATLSX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATLSX0P5H7R 0 0 ;
  SIZE 5.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.8 1.48 ;
        RECT 5.215 1.015 5.305 1.48 ;
        RECT 4.177 1.24 4.317 1.48 ;
        RECT 2.953 1.085 3.043 1.48 ;
        RECT 0.644 1.095 0.784 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.8 0.08 ;
        RECT 5.114 -0.08 5.254 0.16 ;
        RECT 4.064 -0.08 4.204 0.16 ;
        RECT 2.42 -0.08 2.56 0.275 ;
        RECT 0.79 -0.08 0.93 0.26 ;
        RECT 0.32 -0.08 0.41 0.345 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.53 1.35 0.84 ;
        RECT 0.69 0.53 1.35 0.62 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.765 0.425 3.945 0.575 ;
      LAYER MET2 ;
        RECT 3.85 0.23 3.95 0.76 ;
      LAYER VIA1 ;
        RECT 3.855 0.455 3.945 0.545 ;
    END
  END GN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.805 0.88 4.945 0.97 ;
        RECT 4.855 0.363 4.945 0.97 ;
        RECT 4.777 0.35 4.919 0.44 ;
      LAYER MET2 ;
        RECT 4.85 0.23 4.95 0.76 ;
      LAYER VIA1 ;
        RECT 4.855 0.455 4.945 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.455 0.88 4.6 0.97 ;
        RECT 4.455 0.35 4.595 0.44 ;
        RECT 4.455 0.35 4.545 0.97 ;
      LAYER MET2 ;
        RECT 4.45 0.425 4.55 0.96 ;
      LAYER VIA1 ;
        RECT 4.455 0.655 4.545 0.745 ;
    END
  END QN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.57 0.37 0.795 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 3.43 0.96 3.944 1.05 ;
      RECT 5.469 0.25 5.559 1.01 ;
      RECT 2.295 0.7 3.132 0.79 ;
      RECT 2.295 0.57 2.385 0.79 ;
      RECT 5.076 0.25 5.559 0.34 ;
      RECT 4.407 0.17 4.958 0.26 ;
      RECT 5.038 0.231 5.076 0.34 ;
      RECT 4.996 0.191 5.038 0.319 ;
      RECT 4.958 0.17 4.996 0.279 ;
      RECT 4.369 0.17 4.407 0.279 ;
      RECT 4.351 0.179 4.369 0.307 ;
      RECT 4.305 0.211 4.351 0.339 ;
      RECT 4.261 0.256 4.305 0.749 ;
      RECT 4.215 0.301 4.261 0.794 ;
      RECT 4.212 0.69 4.215 0.819 ;
      RECT 4.166 0.715 4.212 0.843 ;
      RECT 4.12 0.761 4.166 0.889 ;
      RECT 4.074 0.807 4.12 0.935 ;
      RECT 4.028 0.853 4.074 0.981 ;
      RECT 3.982 0.899 4.028 1.027 ;
      RECT 3.944 0.941 3.982 1.05 ;
      RECT 3.392 0.941 3.43 1.05 ;
      RECT 3.354 0.903 3.392 1.031 ;
      RECT 3.308 0.861 3.354 0.989 ;
      RECT 3.262 0.815 3.308 0.943 ;
      RECT 3.216 0.769 3.262 0.897 ;
      RECT 3.17 0.723 3.216 0.851 ;
      RECT 3.132 0.7 3.17 0.809 ;
      RECT 3.316 1.14 4.058 1.23 ;
      RECT 3.278 1.083 3.316 1.211 ;
      RECT 3.278 1.14 4.1 1.209 ;
      RECT 3.232 1.14 4.138 1.169 ;
      RECT 5.035 0.685 5.125 1.15 ;
      RECT 4.02 1.121 5.125 1.15 ;
      RECT 4.1 1.06 5.125 1.15 ;
      RECT 3.232 1.121 3.354 1.169 ;
      RECT 3.186 0.995 3.232 1.123 ;
      RECT 4.058 1.081 5.125 1.15 ;
      RECT 3.232 1.041 3.278 1.169 ;
      RECT 3.14 0.949 3.186 1.077 ;
      RECT 3.094 0.903 3.14 1.031 ;
      RECT 3.056 0.949 3.186 0.989 ;
      RECT 1.9 0.88 2.04 0.985 ;
      RECT 1.645 0.88 3.094 0.97 ;
      RECT 1.645 0.17 1.735 0.97 ;
      RECT 1.07 0.17 1.735 0.26 ;
      RECT 3.728 0.78 3.906 0.87 ;
      RECT 3.728 0.78 3.952 0.847 ;
      RECT 3.868 0.761 3.998 0.801 ;
      RECT 3.906 0.719 3.998 0.801 ;
      RECT 3.952 0.673 4.035 0.76 ;
      RECT 4.035 0.282 4.081 0.718 ;
      RECT 4.035 0.327 4.125 0.673 ;
      RECT 3.998 0.631 4.125 0.673 ;
      RECT 4.021 0.252 4.035 0.38 ;
      RECT 3.983 0.327 4.125 0.354 ;
      RECT 3.173 0.245 4.021 0.335 ;
      RECT 3.468 0.78 3.608 0.87 ;
      RECT 3.468 0.52 3.558 0.87 ;
      RECT 1.825 0.365 1.915 0.735 ;
      RECT 2.775 0.52 3.558 0.61 ;
      RECT 2.775 0.315 2.865 0.61 ;
      RECT 1.825 0.365 2.865 0.455 ;
      RECT 0.945 1.1 2.829 1.19 ;
      RECT 2.689 1.06 2.829 1.19 ;
      RECT 0.945 0.725 1.035 1.19 ;
      RECT 0.07 0.255 0.16 1.065 ;
      RECT 0.07 0.915 1.035 1.005 ;
      RECT 0.945 0.725 1.085 0.815 ;
      RECT 1.465 0.35 1.555 1.01 ;
      RECT 0.55 0.35 1.555 0.44 ;
      RECT 0.55 0.275 0.64 0.44 ;
  END
END LATLSX0P5H7R

MACRO LATLSX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATLSX1H7R 0 0 ;
  SIZE 5.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.8 1.48 ;
        RECT 5.215 1.07 5.305 1.48 ;
        RECT 4.177 1.24 4.317 1.48 ;
        RECT 2.953 1.085 3.043 1.48 ;
        RECT 0.644 1.095 0.784 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.8 0.08 ;
        RECT 5.114 -0.08 5.254 0.16 ;
        RECT 4.064 -0.08 4.204 0.16 ;
        RECT 2.42 -0.08 2.56 0.275 ;
        RECT 0.79 -0.08 0.93 0.26 ;
        RECT 0.32 -0.08 0.41 0.345 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.53 1.35 0.84 ;
        RECT 0.69 0.53 1.35 0.62 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.765 0.425 3.945 0.575 ;
      LAYER MET2 ;
        RECT 3.85 0.23 3.95 0.76 ;
      LAYER VIA1 ;
        RECT 3.855 0.455 3.945 0.545 ;
    END
  END GN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.805 0.875 4.945 0.965 ;
        RECT 4.855 0.363 4.945 0.965 ;
        RECT 4.777 0.35 4.919 0.44 ;
      LAYER MET2 ;
        RECT 4.85 0.23 4.95 0.76 ;
      LAYER VIA1 ;
        RECT 4.855 0.455 4.945 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.455 0.87 4.6 0.96 ;
        RECT 4.455 0.35 4.595 0.44 ;
        RECT 4.455 0.35 4.545 0.96 ;
      LAYER MET2 ;
        RECT 4.45 0.425 4.55 0.96 ;
      LAYER VIA1 ;
        RECT 4.455 0.655 4.545 0.745 ;
    END
  END QN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.57 0.37 0.795 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 5.469 0.25 5.559 1.065 ;
      RECT 3.43 0.96 3.944 1.05 ;
      RECT 2.295 0.7 3.132 0.79 ;
      RECT 2.295 0.57 2.385 0.79 ;
      RECT 5.076 0.25 5.559 0.34 ;
      RECT 4.407 0.17 4.958 0.26 ;
      RECT 5.038 0.231 5.076 0.34 ;
      RECT 4.996 0.191 5.038 0.319 ;
      RECT 4.958 0.17 4.996 0.279 ;
      RECT 4.369 0.17 4.407 0.279 ;
      RECT 4.351 0.179 4.369 0.307 ;
      RECT 4.305 0.211 4.351 0.339 ;
      RECT 4.261 0.256 4.305 0.749 ;
      RECT 4.215 0.301 4.261 0.794 ;
      RECT 4.212 0.69 4.215 0.819 ;
      RECT 4.166 0.715 4.212 0.843 ;
      RECT 4.12 0.761 4.166 0.889 ;
      RECT 4.074 0.807 4.12 0.935 ;
      RECT 4.028 0.853 4.074 0.981 ;
      RECT 3.982 0.899 4.028 1.027 ;
      RECT 3.944 0.941 3.982 1.05 ;
      RECT 3.392 0.941 3.43 1.05 ;
      RECT 3.354 0.903 3.392 1.031 ;
      RECT 3.308 0.861 3.354 0.989 ;
      RECT 3.262 0.815 3.308 0.943 ;
      RECT 3.216 0.769 3.262 0.897 ;
      RECT 3.17 0.723 3.216 0.851 ;
      RECT 3.132 0.7 3.17 0.809 ;
      RECT 3.316 1.14 4.058 1.23 ;
      RECT 3.278 1.083 3.316 1.211 ;
      RECT 3.278 1.14 4.1 1.209 ;
      RECT 3.232 1.14 4.138 1.169 ;
      RECT 5.035 0.62 5.125 1.15 ;
      RECT 4.02 1.121 5.125 1.15 ;
      RECT 4.1 1.06 5.125 1.15 ;
      RECT 3.232 1.121 3.354 1.169 ;
      RECT 3.186 0.995 3.232 1.123 ;
      RECT 4.058 1.081 5.125 1.15 ;
      RECT 3.232 1.041 3.278 1.169 ;
      RECT 3.14 0.949 3.186 1.077 ;
      RECT 3.094 0.903 3.14 1.031 ;
      RECT 3.056 0.949 3.186 0.989 ;
      RECT 1.9 0.88 2.04 0.985 ;
      RECT 1.645 0.88 3.094 0.97 ;
      RECT 1.645 0.17 1.735 0.97 ;
      RECT 1.07 0.17 1.735 0.26 ;
      RECT 3.728 0.78 3.906 0.87 ;
      RECT 3.728 0.78 3.952 0.847 ;
      RECT 3.868 0.761 3.998 0.801 ;
      RECT 3.906 0.719 3.998 0.801 ;
      RECT 3.952 0.673 4.035 0.76 ;
      RECT 4.035 0.282 4.081 0.718 ;
      RECT 4.035 0.327 4.125 0.673 ;
      RECT 3.998 0.631 4.125 0.673 ;
      RECT 4.021 0.252 4.035 0.38 ;
      RECT 3.983 0.327 4.125 0.354 ;
      RECT 3.173 0.245 4.021 0.335 ;
      RECT 3.468 0.78 3.608 0.87 ;
      RECT 3.468 0.52 3.558 0.87 ;
      RECT 1.825 0.365 1.915 0.735 ;
      RECT 2.775 0.52 3.558 0.61 ;
      RECT 2.775 0.315 2.865 0.61 ;
      RECT 1.825 0.365 2.865 0.455 ;
      RECT 0.945 1.1 2.829 1.19 ;
      RECT 2.689 1.06 2.829 1.19 ;
      RECT 0.945 0.725 1.035 1.19 ;
      RECT 0.07 0.255 0.16 1.065 ;
      RECT 0.07 0.915 1.035 1.005 ;
      RECT 0.945 0.725 1.085 0.815 ;
      RECT 1.465 0.35 1.555 1.01 ;
      RECT 0.55 0.35 1.555 0.44 ;
      RECT 0.55 0.275 0.64 0.44 ;
  END
END LATLSX1H7R

MACRO LATLSX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATLSX2H7R 0 0 ;
  SIZE 5.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.8 1.48 ;
        RECT 5.215 1.07 5.305 1.48 ;
        RECT 4.177 1.24 4.317 1.48 ;
        RECT 2.953 1.085 3.043 1.48 ;
        RECT 0.644 1.095 0.784 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.8 0.08 ;
        RECT 5.114 -0.08 5.254 0.16 ;
        RECT 4.064 -0.08 4.204 0.16 ;
        RECT 2.42 -0.08 2.56 0.275 ;
        RECT 0.79 -0.08 0.93 0.26 ;
        RECT 0.32 -0.08 0.41 0.345 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.53 1.35 0.84 ;
        RECT 0.69 0.53 1.35 0.62 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.765 0.425 3.945 0.575 ;
      LAYER MET2 ;
        RECT 3.85 0.23 3.95 0.76 ;
      LAYER VIA1 ;
        RECT 3.855 0.455 3.945 0.545 ;
    END
  END GN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.777 0.83 4.945 0.92 ;
        RECT 4.855 0.375 4.945 0.92 ;
        RECT 4.777 0.375 4.945 0.465 ;
      LAYER MET2 ;
        RECT 4.85 0.23 4.95 0.76 ;
      LAYER VIA1 ;
        RECT 4.855 0.455 4.945 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.455 0.83 4.65 0.92 ;
        RECT 4.455 0.375 4.595 0.465 ;
        RECT 4.455 0.375 4.545 0.92 ;
      LAYER MET2 ;
        RECT 4.45 0.425 4.55 0.96 ;
      LAYER VIA1 ;
        RECT 4.455 0.655 4.545 0.745 ;
    END
  END QN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.57 0.37 0.795 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 5.469 0.25 5.559 1.065 ;
      RECT 3.43 0.96 3.944 1.05 ;
      RECT 2.295 0.7 3.132 0.79 ;
      RECT 2.295 0.57 2.385 0.79 ;
      RECT 5.076 0.25 5.559 0.34 ;
      RECT 4.432 0.17 4.958 0.26 ;
      RECT 5.038 0.231 5.076 0.34 ;
      RECT 4.996 0.191 5.038 0.319 ;
      RECT 4.958 0.17 4.996 0.279 ;
      RECT 4.394 0.17 4.432 0.279 ;
      RECT 4.351 0.191 4.394 0.32 ;
      RECT 4.305 0.236 4.351 0.364 ;
      RECT 4.261 0.281 4.305 0.749 ;
      RECT 4.215 0.326 4.261 0.794 ;
      RECT 4.212 0.69 4.215 0.819 ;
      RECT 4.166 0.715 4.212 0.843 ;
      RECT 4.12 0.761 4.166 0.889 ;
      RECT 4.074 0.807 4.12 0.935 ;
      RECT 4.028 0.853 4.074 0.981 ;
      RECT 3.982 0.899 4.028 1.027 ;
      RECT 3.944 0.941 3.982 1.05 ;
      RECT 3.392 0.941 3.43 1.05 ;
      RECT 3.354 0.903 3.392 1.031 ;
      RECT 3.308 0.861 3.354 0.989 ;
      RECT 3.262 0.815 3.308 0.943 ;
      RECT 3.216 0.769 3.262 0.897 ;
      RECT 3.17 0.723 3.216 0.851 ;
      RECT 3.132 0.7 3.17 0.809 ;
      RECT 3.316 1.14 4.058 1.23 ;
      RECT 3.278 1.083 3.316 1.211 ;
      RECT 3.278 1.14 4.1 1.209 ;
      RECT 3.232 1.14 4.138 1.169 ;
      RECT 5.035 0.62 5.125 1.15 ;
      RECT 4.02 1.121 5.125 1.15 ;
      RECT 4.1 1.06 5.125 1.15 ;
      RECT 3.232 1.121 3.354 1.169 ;
      RECT 3.186 0.995 3.232 1.123 ;
      RECT 4.058 1.081 5.125 1.15 ;
      RECT 3.232 1.041 3.278 1.169 ;
      RECT 3.14 0.949 3.186 1.077 ;
      RECT 3.094 0.903 3.14 1.031 ;
      RECT 3.056 0.949 3.186 0.989 ;
      RECT 1.9 0.88 2.04 0.985 ;
      RECT 1.645 0.88 3.094 0.97 ;
      RECT 1.645 0.17 1.735 0.97 ;
      RECT 1.07 0.17 1.735 0.26 ;
      RECT 3.728 0.78 3.906 0.87 ;
      RECT 3.728 0.78 3.952 0.847 ;
      RECT 3.868 0.761 3.998 0.801 ;
      RECT 3.906 0.719 3.998 0.801 ;
      RECT 3.952 0.673 4.035 0.76 ;
      RECT 4.035 0.282 4.081 0.718 ;
      RECT 4.035 0.327 4.125 0.673 ;
      RECT 3.998 0.631 4.125 0.673 ;
      RECT 4.021 0.252 4.035 0.38 ;
      RECT 3.983 0.327 4.125 0.354 ;
      RECT 3.173 0.245 4.021 0.335 ;
      RECT 3.468 0.78 3.608 0.87 ;
      RECT 3.468 0.52 3.558 0.87 ;
      RECT 1.825 0.365 1.915 0.735 ;
      RECT 2.775 0.52 3.558 0.61 ;
      RECT 2.775 0.315 2.865 0.61 ;
      RECT 1.825 0.365 2.865 0.455 ;
      RECT 0.945 1.1 2.829 1.19 ;
      RECT 2.689 1.06 2.829 1.19 ;
      RECT 0.945 0.725 1.035 1.19 ;
      RECT 0.07 0.255 0.16 1.065 ;
      RECT 0.07 0.915 1.035 1.005 ;
      RECT 0.945 0.725 1.085 0.815 ;
      RECT 1.465 0.35 1.555 1.01 ;
      RECT 0.55 0.35 1.555 0.44 ;
      RECT 0.55 0.275 0.64 0.44 ;
  END
END LATLSX2H7R

MACRO LATLX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATLX0P5H7R 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.8 1.48 ;
        RECT 3.355 0.805 3.445 1.48 ;
        RECT 2.78 1.069 2.87 1.48 ;
        RECT 2.1 1.07 2.19 1.48 ;
        RECT 0.828 1.07 0.918 1.48 ;
        RECT 0.336 1.045 0.426 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.8 0.08 ;
        RECT 3.349 -0.08 3.489 0.175 ;
        RECT 2.676 -0.08 2.816 0.174 ;
        RECT 2.075 -0.08 2.165 0.33 ;
        RECT 0.845 -0.08 0.985 0.16 ;
        RECT 0.32 -0.08 0.46 0.175 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.915 0.65 1.185 0.75 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.505 0.35 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END GN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.045 0.815 3.185 0.975 ;
        RECT 3.045 0.35 3.135 0.975 ;
      LAYER MET2 ;
        RECT 3.05 0.63 3.15 1.16 ;
      LAYER VIA1 ;
        RECT 3.055 0.855 3.145 0.945 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.435 0.225 2.525 0.93 ;
        RECT 2.255 0.225 2.525 0.375 ;
      LAYER MET2 ;
        RECT 2.25 0.18 2.35 0.56 ;
      LAYER VIA1 ;
        RECT 2.255 0.255 2.345 0.345 ;
    END
  END QN
  OBS
    LAYER MET1 ;
      RECT 3.62 0.805 3.73 0.945 ;
      RECT 3.64 0.296 3.73 0.945 ;
      RECT 2.615 0.339 2.705 0.696 ;
      RECT 2.615 0.339 2.838 0.429 ;
      RECT 2.615 0.339 2.884 0.406 ;
      RECT 3.303 0.296 3.73 0.386 ;
      RECT 3.261 0.237 3.303 0.365 ;
      RECT 2.781 0.316 2.93 0.36 ;
      RECT 3.215 0.193 3.261 0.321 ;
      RECT 2.827 0.287 2.95 0.327 ;
      RECT 3.215 0.277 3.341 0.321 ;
      RECT 2.838 0.259 2.996 0.294 ;
      RECT 2.93 0.18 2.95 0.327 ;
      RECT 3.177 0.17 3.215 0.279 ;
      RECT 2.838 0.259 3.007 0.266 ;
      RECT 2.95 0.17 3.215 0.26 ;
      RECT 2.884 0.213 2.93 0.36 ;
      RECT 1.585 1.065 2.01 1.155 ;
      RECT 1.92 0.45 2.01 1.155 ;
      RECT 2.358 1.02 2.611 1.11 ;
      RECT 2.354 0.98 2.358 1.108 ;
      RECT 2.354 1.02 2.657 1.087 ;
      RECT 2.308 0.955 2.354 1.083 ;
      RECT 2.262 0.909 2.308 1.037 ;
      RECT 2.573 1.001 2.703 1.041 ;
      RECT 2.262 1.001 2.396 1.037 ;
      RECT 2.611 0.959 2.703 1.041 ;
      RECT 2.224 0.886 2.262 0.995 ;
      RECT 1.92 0.886 2.262 0.976 ;
      RECT 2.657 0.913 2.749 0.995 ;
      RECT 2.703 0.867 2.795 0.949 ;
      RECT 2.703 0.867 2.841 0.903 ;
      RECT 2.749 0.821 2.865 0.868 ;
      RECT 2.795 0.775 2.911 0.833 ;
      RECT 2.841 0.74 2.865 0.868 ;
      RECT 2.865 0.595 2.955 0.788 ;
      RECT 1.895 0.245 1.985 0.525 ;
      RECT 1.385 0.245 1.985 0.335 ;
      RECT 0.07 0.265 0.16 1.055 ;
      RECT 0.07 0.865 0.442 0.955 ;
      RECT 0.07 0.865 0.488 0.932 ;
      RECT 1.715 0.769 1.83 0.909 ;
      RECT 0.404 0.846 0.51 0.898 ;
      RECT 0.442 0.804 0.556 0.864 ;
      RECT 0.488 0.77 0.51 0.898 ;
      RECT 0.51 0.656 0.6 0.819 ;
      RECT 1.715 0.47 1.805 0.909 ;
      RECT 1.255 0.47 1.395 0.58 ;
      RECT 1.036 0.47 1.805 0.56 ;
      RECT 1.015 0.413 1.036 0.55 ;
      RECT 0.969 0.38 1.015 0.516 ;
      RECT 0.923 0.334 0.969 0.47 ;
      RECT 0.923 0.447 1.082 0.47 ;
      RECT 0.877 0.288 0.923 0.424 ;
      RECT 0.831 0.334 0.969 0.378 ;
      RECT 0.07 0.265 0.877 0.355 ;
      RECT 0.578 0.924 0.668 1.087 ;
      RECT 0.578 0.924 0.69 0.975 ;
      RECT 0.578 0.924 0.709 0.955 ;
      RECT 1.51 0.651 1.6 0.945 ;
      RECT 0.624 0.879 1.6 0.945 ;
      RECT 0.668 0.855 1.6 0.945 ;
      RECT 0.668 0.846 0.78 0.945 ;
      RECT 0.69 0.445 0.78 0.945 ;
      RECT 0.565 0.445 0.78 0.535 ;
  END
END LATLX0P5H7R

MACRO LATLX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATLX1H7R 0 0 ;
  SIZE 4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4 1.48 ;
        RECT 3.355 0.805 3.445 1.48 ;
        RECT 2.815 0.995 2.905 1.48 ;
        RECT 2.07 1.07 2.16 1.48 ;
        RECT 0.81 1.07 0.9 1.48 ;
        RECT 0.33 1.045 0.42 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4 0.08 ;
        RECT 3.37 -0.08 3.51 0.175 ;
        RECT 2.655 -0.08 2.795 0.175 ;
        RECT 2.07 -0.08 2.16 0.33 ;
        RECT 0.83 -0.08 0.97 0.175 ;
        RECT 0.32 -0.08 0.46 0.175 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.905 0.655 1.175 0.755 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.505 0.35 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END GN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.055 0.35 3.155 1.13 ;
      LAYER MET2 ;
        RECT 3.05 0.63 3.15 1.16 ;
      LAYER VIA1 ;
        RECT 3.055 0.855 3.145 0.945 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.405 0.32 2.495 0.93 ;
        RECT 2.255 0.32 2.495 0.41 ;
        RECT 2.255 0.225 2.345 0.41 ;
      LAYER MET2 ;
        RECT 2.25 0.18 2.35 0.56 ;
      LAYER VIA1 ;
        RECT 2.255 0.255 2.345 0.345 ;
    END
  END QN
  OBS
    LAYER MET1 ;
      RECT 3.595 0.83 3.75 0.92 ;
      RECT 3.66 0.296 3.75 0.92 ;
      RECT 2.585 0.492 2.675 0.696 ;
      RECT 2.585 0.492 2.721 0.549 ;
      RECT 2.631 0.447 2.767 0.503 ;
      RECT 2.675 0.402 2.813 0.457 ;
      RECT 2.721 0.356 2.859 0.411 ;
      RECT 3.323 0.296 3.75 0.386 ;
      RECT 3.281 0.237 3.323 0.365 ;
      RECT 2.767 0.31 2.905 0.365 ;
      RECT 3.235 0.193 3.281 0.321 ;
      RECT 2.813 0.264 2.93 0.33 ;
      RECT 3.235 0.277 3.361 0.321 ;
      RECT 2.813 0.264 2.976 0.294 ;
      RECT 3.197 0.17 3.235 0.279 ;
      RECT 2.859 0.218 2.987 0.266 ;
      RECT 2.905 0.182 2.93 0.33 ;
      RECT 2.93 0.17 3.235 0.26 ;
      RECT 1.555 1.065 1.98 1.155 ;
      RECT 1.89 0.245 1.98 1.155 ;
      RECT 2.357 1.049 2.542 1.139 ;
      RECT 2.328 0.996 2.357 1.125 ;
      RECT 2.328 1.049 2.588 1.116 ;
      RECT 2.282 0.959 2.328 1.087 ;
      RECT 2.504 1.03 2.634 1.07 ;
      RECT 2.282 1.03 2.395 1.087 ;
      RECT 2.236 0.913 2.282 1.041 ;
      RECT 2.542 0.988 2.634 1.07 ;
      RECT 2.198 0.89 2.236 0.999 ;
      RECT 2.588 0.942 2.68 1.024 ;
      RECT 1.89 0.89 2.236 0.98 ;
      RECT 2.634 0.896 2.726 0.978 ;
      RECT 2.68 0.85 2.772 0.932 ;
      RECT 2.726 0.804 2.813 0.889 ;
      RECT 2.726 0.804 2.851 0.849 ;
      RECT 2.875 0.595 2.965 0.83 ;
      RECT 2.772 0.76 2.965 0.83 ;
      RECT 2.813 0.74 2.965 0.83 ;
      RECT 1.355 0.245 1.98 0.335 ;
      RECT 0.07 0.265 0.16 1.055 ;
      RECT 0.07 0.865 0.457 0.955 ;
      RECT 0.07 0.865 0.503 0.932 ;
      RECT 1.71 0.449 1.8 0.909 ;
      RECT 0.419 0.846 0.556 0.879 ;
      RECT 0.503 0.777 0.51 0.906 ;
      RECT 0.457 0.804 0.556 0.879 ;
      RECT 0.51 0.656 0.6 0.834 ;
      RECT 1.235 0.449 1.375 0.585 ;
      RECT 1.015 0.449 1.8 0.539 ;
      RECT 0.969 0.38 1.015 0.516 ;
      RECT 0.923 0.334 0.969 0.47 ;
      RECT 0.923 0.426 1.061 0.47 ;
      RECT 0.877 0.288 0.923 0.424 ;
      RECT 0.831 0.334 0.969 0.378 ;
      RECT 0.07 0.265 0.877 0.355 ;
      RECT 0.56 0.957 0.65 1.122 ;
      RECT 0.606 0.912 0.724 0.962 ;
      RECT 0.65 0.87 0.69 0.999 ;
      RECT 0.69 0.855 1.365 0.945 ;
      RECT 1.48 0.715 1.57 0.855 ;
      RECT 1.275 0.765 1.57 0.855 ;
      RECT 0.69 0.445 0.78 0.945 ;
      RECT 0.565 0.445 0.78 0.535 ;
  END
END LATLX1H7R

MACRO LATLX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATLX2H7R 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.8 1.48 ;
        RECT 3.255 0.805 3.345 1.48 ;
        RECT 2.73 1.095 2.87 1.48 ;
        RECT 2.06 1.095 2.2 1.48 ;
        RECT 0.32 1.319 1.154 1.48 ;
        RECT 0.8 1.07 0.89 1.48 ;
        RECT 0.32 1.045 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.8 0.08 ;
        RECT 3.314 -0.08 3.454 0.175 ;
        RECT 2.64 -0.08 2.78 0.174 ;
        RECT 2.03 -0.08 2.12 0.33 ;
        RECT 0.82 -0.08 0.96 0.175 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.905 0.655 1.175 0.755 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.505 0.35 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END GN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.01 1.025 3.145 1.175 ;
        RECT 3.01 0.35 3.1 1.175 ;
      LAYER MET2 ;
        RECT 3.05 0.84 3.15 1.22 ;
      LAYER VIA1 ;
        RECT 3.055 1.055 3.145 1.145 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.42 0.485 2.51 0.93 ;
        RECT 2.255 0.485 2.51 0.575 ;
        RECT 2.255 0.335 2.37 0.575 ;
      LAYER MET2 ;
        RECT 2.25 0.23 2.35 0.76 ;
      LAYER VIA1 ;
        RECT 2.255 0.455 2.345 0.545 ;
    END
  END QN
  OBS
    LAYER MET1 ;
      RECT 3.495 0.83 3.695 0.92 ;
      RECT 3.605 0.31 3.695 0.92 ;
      RECT 2.6 0.265 2.69 0.696 ;
      RECT 3.282 0.31 3.695 0.4 ;
      RECT 3.272 0.267 3.282 0.395 ;
      RECT 3.226 0.239 3.272 0.367 ;
      RECT 2.6 0.265 2.877 0.355 ;
      RECT 3.18 0.193 3.226 0.321 ;
      RECT 3.18 0.291 3.32 0.321 ;
      RECT 2.6 0.265 2.961 0.294 ;
      RECT 3.142 0.17 3.18 0.279 ;
      RECT 2.82 0.242 2.972 0.266 ;
      RECT 2.877 0.189 2.915 0.336 ;
      RECT 2.915 0.17 3.18 0.26 ;
      RECT 2.866 0.213 2.877 0.355 ;
      RECT 1.545 1.065 1.97 1.155 ;
      RECT 1.88 0.589 1.97 1.155 ;
      RECT 2.343 1.02 2.586 1.11 ;
      RECT 2.322 0.971 2.343 1.1 ;
      RECT 2.322 1.02 2.632 1.087 ;
      RECT 2.276 0.938 2.322 1.066 ;
      RECT 2.548 1.001 2.691 1.024 ;
      RECT 2.632 0.925 2.653 1.054 ;
      RECT 2.238 1.001 2.381 1.024 ;
      RECT 2.83 0.595 2.92 1.005 ;
      RECT 1.88 0.915 2.276 1.005 ;
      RECT 2.586 0.959 2.92 1.005 ;
      RECT 2.653 0.915 2.92 1.005 ;
      RECT 1.85 0.245 1.94 0.679 ;
      RECT 1.345 0.245 1.94 0.335 ;
      RECT 0.07 0.265 0.16 1.055 ;
      RECT 1.67 0.835 1.79 0.975 ;
      RECT 0.07 0.865 0.442 0.955 ;
      RECT 0.07 0.865 0.488 0.932 ;
      RECT 0.404 0.846 0.51 0.898 ;
      RECT 0.442 0.804 0.556 0.864 ;
      RECT 0.488 0.77 0.51 0.898 ;
      RECT 1.67 0.449 1.76 0.975 ;
      RECT 0.51 0.656 0.6 0.819 ;
      RECT 1.225 0.449 1.365 0.58 ;
      RECT 1.175 0.449 1.76 0.539 ;
      RECT 1.129 0.38 1.175 0.516 ;
      RECT 1.083 0.334 1.129 0.47 ;
      RECT 1.083 0.426 1.221 0.47 ;
      RECT 1.037 0.288 1.083 0.424 ;
      RECT 0.991 0.334 1.129 0.378 ;
      RECT 0.07 0.265 1.037 0.355 ;
      RECT 0.55 0.952 0.64 1.115 ;
      RECT 0.55 0.952 0.686 0.991 ;
      RECT 0.596 0.907 0.69 0.966 ;
      RECT 0.596 0.907 0.719 0.95 ;
      RECT 1.265 0.735 1.355 0.935 ;
      RECT 0.64 0.862 1.355 0.935 ;
      RECT 0.686 0.845 1.355 0.935 ;
      RECT 0.686 0.837 0.78 0.935 ;
      RECT 0.69 0.445 0.78 0.935 ;
      RECT 1.265 0.735 1.56 0.825 ;
      RECT 1.47 0.685 1.56 0.825 ;
      RECT 0.555 0.445 0.78 0.535 ;
  END
END LATLX2H7R

MACRO LATLX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATLX3H7R 0 0 ;
  SIZE 4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4 1.48 ;
        RECT 3.465 0.95 3.555 1.48 ;
        RECT 2.91 1.07 3 1.48 ;
        RECT 2.19 1.061 2.28 1.48 ;
        RECT 0.828 1.07 0.918 1.48 ;
        RECT 0.336 1.045 0.426 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4 0.08 ;
        RECT 3.475 -0.08 3.615 0.175 ;
        RECT 2.72 -0.08 2.86 0.174 ;
        RECT 2.165 -0.08 2.255 0.33 ;
        RECT 0.895 -0.08 1.035 0.16 ;
        RECT 0.32 -0.08 0.46 0.175 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.96 0.65 1.185 0.77 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.505 0.35 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END GN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.155 0.825 3.345 1.03 ;
        RECT 3.155 0.35 3.245 1.03 ;
      LAYER MET2 ;
        RECT 3.25 0.63 3.35 1.16 ;
      LAYER VIA1 ;
        RECT 3.255 0.855 3.345 0.945 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.55 0.655 2.64 1.042 ;
        RECT 2.415 0.655 2.64 0.745 ;
        RECT 2.415 0.28 2.505 0.745 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END QN
  OBS
    LAYER MET1 ;
      RECT 3.69 0.832 3.855 0.922 ;
      RECT 3.765 0.271 3.855 0.922 ;
      RECT 2.73 0.264 2.82 0.696 ;
      RECT 3.388 0.271 3.855 0.361 ;
      RECT 2.73 0.264 2.958 0.354 ;
      RECT 3.371 0.224 3.388 0.353 ;
      RECT 3.325 0.193 3.371 0.321 ;
      RECT 2.73 0.264 3.041 0.294 ;
      RECT 3.287 0.252 3.426 0.279 ;
      RECT 2.901 0.241 3.052 0.266 ;
      RECT 2.958 0.188 2.995 0.336 ;
      RECT 2.995 0.17 3.325 0.26 ;
      RECT 2.947 0.212 2.958 0.354 ;
      RECT 2.37 1.14 2.82 1.23 ;
      RECT 2.73 0.786 2.82 1.23 ;
      RECT 1.693 1.08 1.945 1.17 ;
      RECT 1.693 1.08 1.991 1.147 ;
      RECT 2.37 0.847 2.46 1.23 ;
      RECT 1.907 1.061 2.037 1.101 ;
      RECT 1.945 1.019 2.05 1.07 ;
      RECT 2.037 0.948 2.04 1.077 ;
      RECT 1.991 0.973 2.096 1.042 ;
      RECT 2.04 0.589 2.13 1.002 ;
      RECT 2.04 0.847 2.176 0.962 ;
      RECT 2.04 0.847 2.178 0.938 ;
      RECT 2.04 0.847 2.46 0.937 ;
      RECT 2.73 0.786 3.065 0.876 ;
      RECT 2.975 0.556 3.065 0.876 ;
      RECT 1.96 0.261 2.05 0.679 ;
      RECT 1.455 0.261 2.05 0.351 ;
      RECT 0.07 0.265 0.16 1.055 ;
      RECT 0.07 0.865 0.467 0.955 ;
      RECT 1.78 0.769 1.95 0.909 ;
      RECT 0.51 0.656 0.556 0.889 ;
      RECT 0.429 0.846 0.556 0.889 ;
      RECT 0.467 0.805 0.51 0.934 ;
      RECT 0.51 0.656 0.6 0.844 ;
      RECT 1.78 0.449 1.87 0.909 ;
      RECT 1.348 0.449 1.438 0.62 ;
      RECT 1.217 0.449 1.87 0.539 ;
      RECT 1.217 0.25 1.307 0.539 ;
      RECT 0.07 0.265 0.537 0.355 ;
      RECT 0.819 0.25 1.307 0.34 ;
      RECT 0.778 0.191 0.819 0.32 ;
      RECT 0.74 0.25 1.307 0.28 ;
      RECT 0.499 0.246 0.631 0.28 ;
      RECT 0.583 0.176 0.593 0.304 ;
      RECT 0.593 0.171 0.778 0.261 ;
      RECT 0.819 0.231 0.857 0.34 ;
      RECT 0.537 0.204 0.583 0.332 ;
      RECT 0.578 0.965 0.668 1.147 ;
      RECT 0.624 0.92 0.73 0.985 ;
      RECT 0.668 0.887 0.69 1.016 ;
      RECT 0.624 0.92 0.745 0.958 ;
      RECT 1.6 0.68 1.69 0.95 ;
      RECT 0.69 0.86 1.69 0.95 ;
      RECT 0.69 0.446 0.78 0.95 ;
      RECT 0.64 0.38 0.73 0.536 ;
  END
END LATLX3H7R

MACRO LATLX4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LATLX4H7R 0 0 ;
  SIZE 4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4 1.48 ;
        RECT 3.435 0.95 3.525 1.48 ;
        RECT 2.91 1.07 3 1.48 ;
        RECT 2.19 1.07 2.28 1.48 ;
        RECT 0.828 1.07 0.918 1.48 ;
        RECT 0.336 1.045 0.426 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4 0.08 ;
        RECT 3.46 -0.08 3.6 0.175 ;
        RECT 2.72 -0.08 2.86 0.174 ;
        RECT 2.165 -0.08 2.255 0.33 ;
        RECT 0.895 -0.08 1.035 0.16 ;
        RECT 0.32 -0.08 0.46 0.175 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.885 0.655 1.185 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.505 0.35 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END GN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.155 0.825 3.345 0.975 ;
        RECT 3.155 0.35 3.245 0.975 ;
      LAYER MET2 ;
        RECT 3.25 0.63 3.35 1.16 ;
      LAYER VIA1 ;
        RECT 3.255 0.855 3.345 0.945 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.55 0.655 2.64 0.93 ;
        RECT 2.415 0.655 2.64 0.745 ;
        RECT 2.415 0.35 2.505 0.745 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END QN
  OBS
    LAYER MET1 ;
      RECT 3.66 0.832 3.84 0.922 ;
      RECT 3.75 0.271 3.84 0.922 ;
      RECT 2.73 0.264 2.82 0.696 ;
      RECT 3.388 0.271 3.84 0.361 ;
      RECT 2.73 0.264 2.958 0.354 ;
      RECT 3.371 0.224 3.388 0.353 ;
      RECT 3.325 0.193 3.371 0.321 ;
      RECT 2.73 0.264 3.041 0.294 ;
      RECT 3.287 0.252 3.426 0.279 ;
      RECT 2.901 0.241 3.052 0.266 ;
      RECT 2.958 0.188 2.995 0.336 ;
      RECT 2.995 0.17 3.325 0.26 ;
      RECT 2.947 0.212 2.958 0.354 ;
      RECT 1.693 1.065 1.96 1.155 ;
      RECT 1.693 1.065 2.006 1.132 ;
      RECT 2.37 1.02 2.82 1.11 ;
      RECT 2.73 0.786 2.82 1.11 ;
      RECT 1.922 1.046 2.04 1.092 ;
      RECT 1.96 1.004 2.075 1.058 ;
      RECT 2.006 0.964 2.04 1.092 ;
      RECT 2.37 0.89 2.46 1.11 ;
      RECT 2.04 0.429 2.121 1.017 ;
      RECT 2.04 0.429 2.13 0.99 ;
      RECT 2.006 0.964 2.135 0.983 ;
      RECT 2.04 0.89 2.46 0.98 ;
      RECT 2.73 0.786 3.065 0.876 ;
      RECT 2.975 0.556 3.065 0.876 ;
      RECT 1.985 0.261 2.075 0.519 ;
      RECT 1.455 0.261 2.075 0.351 ;
      RECT 0.07 0.265 0.16 1.055 ;
      RECT 0.07 0.865 0.432 0.955 ;
      RECT 0.07 0.865 0.478 0.932 ;
      RECT 1.805 0.769 1.95 0.909 ;
      RECT 0.394 0.846 0.51 0.893 ;
      RECT 0.432 0.804 0.556 0.854 ;
      RECT 0.478 0.765 0.51 0.893 ;
      RECT 0.51 0.641 0.6 0.809 ;
      RECT 1.805 0.47 1.895 0.909 ;
      RECT 1.348 0.47 1.438 0.62 ;
      RECT 1.217 0.47 1.895 0.56 ;
      RECT 1.217 0.25 1.307 0.56 ;
      RECT 0.07 0.265 0.537 0.355 ;
      RECT 0.819 0.25 1.307 0.34 ;
      RECT 0.778 0.191 0.819 0.32 ;
      RECT 0.74 0.25 1.307 0.28 ;
      RECT 0.499 0.246 0.631 0.28 ;
      RECT 0.583 0.176 0.593 0.304 ;
      RECT 0.593 0.171 0.778 0.261 ;
      RECT 0.819 0.231 0.857 0.34 ;
      RECT 0.537 0.204 0.583 0.332 ;
      RECT 0.578 0.915 0.668 1.082 ;
      RECT 0.578 0.915 0.69 0.966 ;
      RECT 0.578 0.915 0.72 0.94 ;
      RECT 1.6 0.68 1.69 0.925 ;
      RECT 0.624 0.87 1.69 0.925 ;
      RECT 0.69 0.835 1.69 0.925 ;
      RECT 0.668 0.837 1.69 0.925 ;
      RECT 0.69 0.446 0.78 0.925 ;
      RECT 0.64 0.38 0.73 0.536 ;
  END
END LATLX4H7R

MACRO MDFFQX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MDFFQX0P5H7R 0 0 ;
  SIZE 6.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.4 1.48 ;
        RECT 5.975 1.07 6.065 1.48 ;
        RECT 5.305 1.24 5.445 1.48 ;
        RECT 3.965 1.05 4.055 1.48 ;
        RECT 3.015 1.24 3.155 1.48 ;
        RECT 1.665 1.05 1.755 1.48 ;
        RECT 0.325 1.11 0.465 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.4 0.08 ;
        RECT 5.605 -0.08 5.695 0.33 ;
        RECT 5.045 -0.08 5.135 0.365 ;
        RECT 4.045 -0.08 4.135 0.365 ;
        RECT 2.875 -0.08 3.015 0.16 ;
        RECT 1.435 -0.08 1.575 0.185 ;
        RECT 0.325 -0.08 0.465 0.185 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.655 0.625 1.835 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END CK
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.48 0.455 0.575 0.645 ;
        RECT 0.38 0.455 0.575 0.545 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.35 0.455 1.575 0.575 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END D1
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.615 0.455 5.705 1.005 ;
        RECT 5.355 0.455 5.705 0.545 ;
        RECT 5.355 0.255 5.445 0.545 ;
      LAYER MET2 ;
        RECT 5.45 0.225 5.55 0.76 ;
      LAYER VIA1 ;
        RECT 5.455 0.455 5.545 0.545 ;
    END
  END Q
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.745 0.855 0.835 ;
        RECT 0.225 0.655 0.375 0.835 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END S0
  OBS
    LAYER MET1 ;
      RECT 5 1.14 5.161 1.23 ;
      RECT 5.518 1.095 5.885 1.185 ;
      RECT 5 1.14 5.241 1.169 ;
      RECT 5.483 1.095 5.885 1.168 ;
      RECT 5.203 1.06 5.521 1.15 ;
      RECT 5.123 1.121 5.885 1.15 ;
      RECT 5.161 1.081 5.203 1.209 ;
      RECT 5.795 0.89 5.885 1.185 ;
      RECT 5.518 1.077 5.556 1.185 ;
      RECT 5.795 0.89 6.355 0.98 ;
      RECT 5.855 0.255 5.945 0.98 ;
      RECT 4.47 0.93 5.115 1.02 ;
      RECT 5.025 0.505 5.115 1.02 ;
      RECT 5.025 0.67 5.525 0.76 ;
      RECT 4.815 0.505 5.115 0.595 ;
      RECT 4.815 0.255 4.905 0.595 ;
      RECT 4.48 0.255 4.905 0.345 ;
      RECT 3.605 0.55 3.695 1.05 ;
      RECT 4.845 0.685 4.935 0.835 ;
      RECT 4.635 0.685 4.935 0.775 ;
      RECT 4.635 0.485 4.725 0.775 ;
      RECT 2.485 0.44 2.575 0.655 ;
      RECT 3.685 0.17 3.775 0.64 ;
      RECT 3.685 0.485 4.725 0.575 ;
      RECT 2.485 0.44 2.69 0.53 ;
      RECT 2.6 0.25 2.69 0.53 ;
      RECT 2.6 0.25 3.092 0.34 ;
      RECT 2.6 0.25 3.172 0.279 ;
      RECT 3.134 0.17 3.775 0.26 ;
      RECT 3.054 0.231 3.775 0.26 ;
      RECT 3.092 0.191 3.134 0.319 ;
      RECT 3.273 1.14 3.875 1.23 ;
      RECT 3.785 0.73 3.875 1.23 ;
      RECT 1.925 1.14 2.897 1.23 ;
      RECT 3.231 1.14 3.875 1.209 ;
      RECT 1.925 1.14 2.939 1.209 ;
      RECT 3.193 1.14 3.875 1.169 ;
      RECT 1.925 1.14 2.977 1.169 ;
      RECT 2.939 1.06 3.231 1.15 ;
      RECT 2.859 1.121 3.311 1.15 ;
      RECT 1.925 0.35 2.015 1.23 ;
      RECT 2.897 1.081 3.273 1.15 ;
      RECT 3.785 0.73 4.52 0.82 ;
      RECT 1.85 0.35 2.015 0.44 ;
      RECT 3.345 0.375 3.435 1.045 ;
      RECT 2.86 0.435 2.95 0.625 ;
      RECT 2.86 0.435 3.435 0.525 ;
      RECT 3.2 0.375 3.57 0.465 ;
      RECT 2.51 0.915 2.866 1.005 ;
      RECT 2.51 0.915 2.901 0.988 ;
      RECT 3.09 0.695 3.18 0.97 ;
      RECT 2.828 0.897 3.18 0.97 ;
      RECT 2.863 0.88 3.18 0.97 ;
      RECT 2.51 0.75 2.6 1.005 ;
      RECT 2.3 0.75 2.6 0.84 ;
      RECT 2.3 0.26 2.39 0.84 ;
      RECT 2.3 0.26 2.485 0.35 ;
      RECT 0.945 0.275 1.035 1.03 ;
      RECT 2.12 0.93 2.34 1.02 ;
      RECT 2.12 0.17 2.21 1.02 ;
      RECT 0.945 0.275 1.755 0.365 ;
      RECT 1.665 0.17 1.755 0.365 ;
      RECT 1.665 0.17 2.21 0.26 ;
      RECT 0.765 1.12 1.395 1.21 ;
      RECT 1.305 0.72 1.395 1.21 ;
      RECT 0.765 0.93 0.855 1.21 ;
      RECT 0.045 0.93 0.855 1.02 ;
      RECT 0.045 0.275 0.135 1.02 ;
      RECT 0.74 0.275 0.83 0.6 ;
      RECT 0.045 0.275 0.83 0.365 ;
  END
END MDFFQX0P5H7R

MACRO MDFFQX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MDFFQX1H7R 0 0 ;
  SIZE 6.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.4 1.48 ;
        RECT 5.99 1.07 6.08 1.48 ;
        RECT 5.305 1.24 5.445 1.48 ;
        RECT 3.965 1.05 4.055 1.48 ;
        RECT 3.015 1.24 3.155 1.48 ;
        RECT 1.665 1.05 1.755 1.48 ;
        RECT 0.325 1.11 0.465 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.4 0.08 ;
        RECT 5.605 -0.08 5.695 0.33 ;
        RECT 5.045 -0.08 5.135 0.365 ;
        RECT 4.045 -0.08 4.135 0.365 ;
        RECT 2.875 -0.08 3.015 0.16 ;
        RECT 1.435 -0.08 1.575 0.185 ;
        RECT 0.325 -0.08 0.465 0.185 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.655 0.625 1.835 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END CK
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.48 0.455 0.575 0.645 ;
        RECT 0.38 0.455 0.575 0.545 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.35 0.455 1.575 0.575 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END D1
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.62 0.455 5.71 1.005 ;
        RECT 5.355 0.455 5.71 0.545 ;
        RECT 5.355 0.295 5.445 0.545 ;
      LAYER MET2 ;
        RECT 5.45 0.225 5.55 0.76 ;
      LAYER VIA1 ;
        RECT 5.455 0.455 5.545 0.545 ;
    END
  END Q
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.745 0.855 0.835 ;
        RECT 0.225 0.655 0.375 0.835 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END S0
  OBS
    LAYER MET1 ;
      RECT 5 1.14 5.161 1.23 ;
      RECT 5.518 1.095 5.89 1.185 ;
      RECT 5 1.14 5.241 1.169 ;
      RECT 5.483 1.095 5.89 1.168 ;
      RECT 5.203 1.06 5.521 1.15 ;
      RECT 5.123 1.121 5.89 1.15 ;
      RECT 5.161 1.081 5.203 1.209 ;
      RECT 5.8 0.89 5.89 1.185 ;
      RECT 5.518 1.077 5.556 1.185 ;
      RECT 6.24 0.89 6.33 1.045 ;
      RECT 5.8 0.89 6.33 0.98 ;
      RECT 5.855 0.275 5.945 0.98 ;
      RECT 4.47 0.93 5.115 1.02 ;
      RECT 5.025 0.505 5.115 1.02 ;
      RECT 5.025 0.67 5.53 0.76 ;
      RECT 4.815 0.505 5.115 0.595 ;
      RECT 4.815 0.255 4.905 0.595 ;
      RECT 4.48 0.255 4.905 0.345 ;
      RECT 3.605 0.55 3.695 1.05 ;
      RECT 4.845 0.685 4.935 0.835 ;
      RECT 4.635 0.685 4.935 0.775 ;
      RECT 4.635 0.485 4.725 0.775 ;
      RECT 2.485 0.44 2.575 0.655 ;
      RECT 3.685 0.17 3.775 0.64 ;
      RECT 3.685 0.485 4.725 0.575 ;
      RECT 2.485 0.44 2.69 0.53 ;
      RECT 2.6 0.25 2.69 0.53 ;
      RECT 2.6 0.25 3.092 0.34 ;
      RECT 2.6 0.25 3.172 0.279 ;
      RECT 3.134 0.17 3.775 0.26 ;
      RECT 3.054 0.231 3.775 0.26 ;
      RECT 3.092 0.191 3.134 0.319 ;
      RECT 3.273 1.14 3.875 1.23 ;
      RECT 3.785 0.73 3.875 1.23 ;
      RECT 1.925 1.14 2.897 1.23 ;
      RECT 3.231 1.14 3.875 1.209 ;
      RECT 1.925 1.14 2.939 1.209 ;
      RECT 3.193 1.14 3.875 1.169 ;
      RECT 1.925 1.14 2.977 1.169 ;
      RECT 2.939 1.06 3.231 1.15 ;
      RECT 2.859 1.121 3.311 1.15 ;
      RECT 1.925 0.35 2.015 1.23 ;
      RECT 2.897 1.081 3.273 1.15 ;
      RECT 3.785 0.73 4.52 0.82 ;
      RECT 1.85 0.35 2.015 0.44 ;
      RECT 3.345 0.375 3.435 1.045 ;
      RECT 2.86 0.435 2.95 0.625 ;
      RECT 2.86 0.435 3.435 0.525 ;
      RECT 3.2 0.375 3.57 0.465 ;
      RECT 2.51 0.915 2.866 1.005 ;
      RECT 2.51 0.915 2.901 0.988 ;
      RECT 3.09 0.695 3.18 0.97 ;
      RECT 2.828 0.897 3.18 0.97 ;
      RECT 2.863 0.88 3.18 0.97 ;
      RECT 2.51 0.75 2.6 1.005 ;
      RECT 2.3 0.75 2.6 0.84 ;
      RECT 2.3 0.26 2.39 0.84 ;
      RECT 2.3 0.26 2.485 0.35 ;
      RECT 0.945 0.275 1.035 1.03 ;
      RECT 2.12 0.93 2.34 1.02 ;
      RECT 2.12 0.17 2.21 1.02 ;
      RECT 0.945 0.275 1.755 0.365 ;
      RECT 1.665 0.17 1.755 0.365 ;
      RECT 1.665 0.17 2.21 0.26 ;
      RECT 0.765 1.12 1.395 1.21 ;
      RECT 1.305 0.72 1.395 1.21 ;
      RECT 0.765 0.93 0.855 1.21 ;
      RECT 0.045 0.93 0.855 1.02 ;
      RECT 0.045 0.275 0.135 1.02 ;
      RECT 0.74 0.275 0.83 0.6 ;
      RECT 0.045 0.275 0.83 0.365 ;
  END
END MDFFQX1H7R

MACRO MDFFQX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MDFFQX2H7R 0 0 ;
  SIZE 6.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.4 1.48 ;
        RECT 5.99 1.07 6.08 1.48 ;
        RECT 5.305 1.24 5.445 1.48 ;
        RECT 3.965 1.05 4.055 1.48 ;
        RECT 3.015 1.24 3.155 1.48 ;
        RECT 1.665 1.05 1.755 1.48 ;
        RECT 0.325 1.11 0.465 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.4 0.08 ;
        RECT 5.605 -0.08 5.695 0.35 ;
        RECT 5.045 -0.08 5.135 0.365 ;
        RECT 4.045 -0.08 4.135 0.365 ;
        RECT 2.875 -0.08 3.015 0.16 ;
        RECT 1.435 -0.08 1.575 0.185 ;
        RECT 0.325 -0.08 0.465 0.185 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.655 0.625 1.835 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END CK
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.48 0.455 0.575 0.645 ;
        RECT 0.38 0.455 0.575 0.545 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.35 0.455 1.575 0.575 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END D1
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.62 0.455 5.71 1.03 ;
        RECT 5.355 0.455 5.71 0.545 ;
        RECT 5.355 0.225 5.445 0.545 ;
      LAYER MET2 ;
        RECT 5.45 0.225 5.55 0.76 ;
      LAYER VIA1 ;
        RECT 5.455 0.455 5.545 0.545 ;
    END
  END Q
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.745 0.855 0.835 ;
        RECT 0.225 0.655 0.375 0.835 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END S0
  OBS
    LAYER MET1 ;
      RECT 5.563 1.14 5.89 1.23 ;
      RECT 5 1.14 5.161 1.23 ;
      RECT 5.521 1.14 5.89 1.209 ;
      RECT 5 1.14 5.203 1.209 ;
      RECT 5.483 1.14 5.89 1.169 ;
      RECT 5 1.14 5.241 1.169 ;
      RECT 5.203 1.06 5.521 1.15 ;
      RECT 5.8 0.89 5.89 1.23 ;
      RECT 5.123 1.121 5.601 1.15 ;
      RECT 5.161 1.081 5.563 1.15 ;
      RECT 5.8 0.89 6.355 0.98 ;
      RECT 5.855 0.31 5.945 0.98 ;
      RECT 4.47 0.93 5.115 1.02 ;
      RECT 5.025 0.505 5.115 1.02 ;
      RECT 5.025 0.67 5.47 0.76 ;
      RECT 4.815 0.505 5.115 0.595 ;
      RECT 4.815 0.255 4.905 0.595 ;
      RECT 4.48 0.255 4.905 0.345 ;
      RECT 3.605 0.55 3.695 1.05 ;
      RECT 4.845 0.685 4.935 0.835 ;
      RECT 4.635 0.685 4.935 0.775 ;
      RECT 4.635 0.485 4.725 0.775 ;
      RECT 2.485 0.44 2.575 0.655 ;
      RECT 3.685 0.17 3.775 0.64 ;
      RECT 3.685 0.485 4.725 0.575 ;
      RECT 2.485 0.44 2.69 0.53 ;
      RECT 2.6 0.25 2.69 0.53 ;
      RECT 2.6 0.25 3.092 0.34 ;
      RECT 2.6 0.25 3.172 0.279 ;
      RECT 3.134 0.17 3.775 0.26 ;
      RECT 3.054 0.231 3.775 0.26 ;
      RECT 3.092 0.191 3.134 0.319 ;
      RECT 3.273 1.14 3.875 1.23 ;
      RECT 3.785 0.73 3.875 1.23 ;
      RECT 1.925 1.14 2.897 1.23 ;
      RECT 3.231 1.14 3.875 1.209 ;
      RECT 1.925 1.14 2.939 1.209 ;
      RECT 3.193 1.14 3.875 1.169 ;
      RECT 1.925 1.14 2.977 1.169 ;
      RECT 2.939 1.06 3.231 1.15 ;
      RECT 2.859 1.121 3.311 1.15 ;
      RECT 1.925 0.35 2.015 1.23 ;
      RECT 2.897 1.081 3.273 1.15 ;
      RECT 3.785 0.73 4.52 0.82 ;
      RECT 1.85 0.35 2.015 0.44 ;
      RECT 3.345 0.375 3.435 1.045 ;
      RECT 2.86 0.435 2.95 0.625 ;
      RECT 2.86 0.435 3.435 0.525 ;
      RECT 3.2 0.375 3.57 0.465 ;
      RECT 2.51 0.915 2.866 1.005 ;
      RECT 2.51 0.915 2.901 0.988 ;
      RECT 3.09 0.695 3.18 0.97 ;
      RECT 2.828 0.897 3.18 0.97 ;
      RECT 2.863 0.88 3.18 0.97 ;
      RECT 2.51 0.75 2.6 1.005 ;
      RECT 2.3 0.75 2.6 0.84 ;
      RECT 2.3 0.26 2.39 0.84 ;
      RECT 2.3 0.26 2.485 0.35 ;
      RECT 0.945 0.275 1.035 1.03 ;
      RECT 2.12 0.93 2.34 1.02 ;
      RECT 2.12 0.17 2.21 1.02 ;
      RECT 0.945 0.275 1.755 0.365 ;
      RECT 1.665 0.17 1.755 0.365 ;
      RECT 1.665 0.17 2.21 0.26 ;
      RECT 0.765 1.12 1.395 1.21 ;
      RECT 1.305 0.72 1.395 1.21 ;
      RECT 0.765 0.93 0.855 1.21 ;
      RECT 0.045 0.93 0.855 1.02 ;
      RECT 0.045 0.275 0.135 1.02 ;
      RECT 0.74 0.275 0.83 0.6 ;
      RECT 0.045 0.275 0.83 0.365 ;
  END
END MDFFQX2H7R

MACRO MSDFFQX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MSDFFQX0P5H7R 0 0 ;
  SIZE 7.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7.4 1.48 ;
        RECT 6.906 0.925 6.996 1.48 ;
        RECT 6.417 1.19 6.557 1.48 ;
        RECT 5.707 1.225 5.852 1.48 ;
        RECT 4.657 1.225 4.797 1.48 ;
        RECT 3.508 1.225 3.648 1.48 ;
        RECT 2.593 1.225 2.733 1.48 ;
        RECT 1.478 1.24 1.618 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7.4 0.08 ;
        RECT 6.922 -0.08 7.012 0.385 ;
        RECT 6.427 -0.08 6.517 0.425 ;
        RECT 5.712 -0.08 5.852 0.175 ;
        RECT 4.567 -0.08 4.707 0.175 ;
        RECT 3.548 -0.08 3.638 0.33 ;
        RECT 2.482 -0.08 2.622 0.175 ;
        RECT 1.525 -0.08 1.615 0.201 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.365 0.625 3.545 0.775 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END CK
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.455 0.575 0.65 ;
        RECT 0.415 0.455 0.575 0.545 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.254 0.705 1.354 0.975 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END D1
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.172 0.625 7.345 0.775 ;
        RECT 7.172 0.31 7.262 0.925 ;
      LAYER MET2 ;
        RECT 7.25 0.425 7.35 0.96 ;
      LAYER VIA1 ;
        RECT 7.255 0.655 7.345 0.745 ;
    END
  END Q
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.925 0.505 1.265 0.595 ;
        RECT 0.225 0.765 1.015 0.855 ;
        RECT 0.925 0.505 1.015 0.855 ;
        RECT 0.225 0.625 0.345 0.855 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END S0
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.763 0.55 2.853 0.714 ;
        RECT 2.688 0.505 2.809 0.554 ;
        RECT 2.21 0.463 2.763 0.535 ;
        RECT 2.726 0.55 2.853 0.592 ;
        RECT 2.21 0.456 2.726 0.535 ;
        RECT 2.233 0.445 2.726 0.535 ;
        RECT 2.118 0.537 2.233 0.585 ;
        RECT 2.164 0.491 2.271 0.554 ;
        RECT 2.072 0.583 2.21 0.619 ;
        RECT 2.023 0.653 2.164 0.665 ;
        RECT 2.026 0.629 2.164 0.665 ;
        RECT 2.072 0.583 2.164 0.665 ;
        RECT 1.825 0.655 2.118 0.711 ;
        RECT 1.825 0.655 2.072 0.757 ;
        RECT 1.825 0.655 2.026 0.78 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.453 0.625 2.633 0.775 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.967 0.96 6.057 1.175 ;
      RECT 5.967 1.01 6.816 1.1 ;
      RECT 6.726 0.745 6.816 1.1 ;
      RECT 5.197 0.96 6.195 1.05 ;
      RECT 6.105 0.31 6.195 1.1 ;
      RECT 5.197 0.35 5.287 1.05 ;
      RECT 6.726 0.745 6.984 0.835 ;
      RECT 6.894 0.559 6.984 0.835 ;
      RECT 5.177 0.35 5.317 0.44 ;
      RECT 5.942 0.31 6.195 0.4 ;
      RECT 6.546 0.565 6.636 0.92 ;
      RECT 6.332 0.565 6.747 0.655 ;
      RECT 6.657 0.287 6.747 0.655 ;
      RECT 5.417 0.78 5.557 0.87 ;
      RECT 5.447 0.7 5.918 0.79 ;
      RECT 5.447 0.17 5.537 0.87 ;
      RECT 5.392 0.512 5.537 0.652 ;
      RECT 4.461 0.27 4.789 0.36 ;
      RECT 4.445 0.224 4.461 0.352 ;
      RECT 4.445 0.27 4.835 0.337 ;
      RECT 4.399 0.193 4.445 0.321 ;
      RECT 4.751 0.251 4.889 0.279 ;
      RECT 4.835 0.178 4.851 0.306 ;
      RECT 4.361 0.251 4.499 0.279 ;
      RECT 4.851 0.17 5.537 0.26 ;
      RECT 4.192 0.17 4.399 0.26 ;
      RECT 4.789 0.209 5.537 0.26 ;
      RECT 4.931 1.14 5.442 1.23 ;
      RECT 3.832 1.14 4.392 1.23 ;
      RECT 4.302 1.045 4.392 1.23 ;
      RECT 4.92 1.096 4.931 1.225 ;
      RECT 4.874 1.068 4.92 1.196 ;
      RECT 3.243 1.075 3.428 1.165 ;
      RECT 4.836 1.121 4.969 1.154 ;
      RECT 3.832 0.42 3.922 1.23 ;
      RECT 4.302 1.045 4.874 1.135 ;
      RECT 3.338 1.045 3.922 1.135 ;
      RECT 3.832 0.522 4.027 0.612 ;
      RECT 3.303 0.42 3.922 0.51 ;
      RECT 3.303 0.205 3.393 0.51 ;
      RECT 3.298 0.205 3.393 0.345 ;
      RECT 4.922 0.865 5.086 0.96 ;
      RECT 4.996 0.35 5.086 0.96 ;
      RECT 4.567 0.865 5.086 0.955 ;
      RECT 4.567 0.678 4.657 0.955 ;
      RECT 4.927 0.35 5.086 0.44 ;
      RECT 4.026 0.847 4.207 0.987 ;
      RECT 4.117 0.422 4.207 0.987 ;
      RECT 4.797 0.543 4.887 0.71 ;
      RECT 4.778 0.543 4.887 0.585 ;
      RECT 4.117 0.485 4.816 0.575 ;
      RECT 4.117 0.508 4.862 0.575 ;
      RECT 4.117 0.464 4.248 0.575 ;
      RECT 4.102 0.346 4.117 0.475 ;
      RECT 4.058 0.377 4.163 0.445 ;
      RECT 4.012 0.228 4.102 0.4 ;
      RECT 2.069 1.05 2.54 1.14 ;
      RECT 2.069 1.05 2.545 1.138 ;
      RECT 2.069 1.05 3.032 1.135 ;
      RECT 2.069 1.05 3.078 1.112 ;
      RECT 2.502 1.047 3.123 1.067 ;
      RECT 2.507 1.045 3.123 1.067 ;
      RECT 2.994 1.026 3.123 1.067 ;
      RECT 3.032 0.984 3.123 1.067 ;
      RECT 3.032 0.984 3.169 1.021 ;
      RECT 3.078 0.938 3.172 0.997 ;
      RECT 3.123 0.392 3.212 0.975 ;
      RECT 3.652 0.6 3.742 0.955 ;
      RECT 3.123 0.865 3.742 0.955 ;
      RECT 3.123 0.412 3.213 0.955 ;
      RECT 3.082 0.171 3.172 0.431 ;
      RECT 1.95 0.265 2.699 0.355 ;
      RECT 1.95 0.265 2.745 0.332 ;
      RECT 2.661 0.246 2.793 0.28 ;
      RECT 2.745 0.176 2.755 0.304 ;
      RECT 2.755 0.171 3.172 0.261 ;
      RECT 2.699 0.204 3.172 0.261 ;
      RECT 1.628 0.87 2.363 0.96 ;
      RECT 2.273 0.685 2.363 0.96 ;
      RECT 1.628 0.87 2.954 0.955 ;
      RECT 1.628 0.87 2.992 0.936 ;
      RECT 2.943 0.468 3.033 0.897 ;
      RECT 2.273 0.865 3.033 0.897 ;
      RECT 2.858 0.809 2.954 0.955 ;
      RECT 1.628 0.549 1.718 0.96 ;
      RECT 2.902 0.351 2.992 0.507 ;
      RECT 2.852 0.351 2.992 0.441 ;
      RECT 0.765 1.065 1.423 1.155 ;
      RECT 1.388 1.06 1.959 1.15 ;
      RECT 1.444 0.3 1.534 1.15 ;
      RECT 0.943 0.3 1.84 0.39 ;
      RECT 0.045 0.925 0.16 1.065 ;
      RECT 0.045 0.27 0.135 1.065 ;
      RECT 0.745 0.27 0.835 0.62 ;
      RECT 0.045 0.27 0.835 0.36 ;
  END
END MSDFFQX0P5H7R

MACRO MSDFFQX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MSDFFQX1H7R 0 0 ;
  SIZE 7.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7.4 1.48 ;
        RECT 6.906 0.93 6.996 1.48 ;
        RECT 6.441 1.23 6.581 1.48 ;
        RECT 5.707 1.225 5.852 1.48 ;
        RECT 4.657 1.225 4.797 1.48 ;
        RECT 3.508 1.225 3.648 1.48 ;
        RECT 2.593 1.225 2.733 1.48 ;
        RECT 1.478 1.24 1.618 1.48 ;
        RECT 0.304 1.092 0.444 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7.4 0.08 ;
        RECT 6.922 -0.08 7.012 0.469 ;
        RECT 6.427 -0.08 6.517 0.425 ;
        RECT 5.712 -0.08 5.852 0.175 ;
        RECT 4.555 -0.08 4.707 0.175 ;
        RECT 3.548 -0.08 3.638 0.33 ;
        RECT 2.482 -0.08 2.622 0.175 ;
        RECT 1.563 -0.08 1.653 0.201 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.303 0.6 3.562 0.775 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END CK
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.455 0.609 0.645 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.178 0.844 1.38 0.97 ;
        RECT 1.221 0.71 1.38 0.97 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END D1
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.172 0.26 7.345 0.945 ;
      LAYER MET2 ;
        RECT 7.25 0.425 7.35 0.96 ;
      LAYER VIA1 ;
        RECT 7.255 0.655 7.345 0.745 ;
    END
  END Q
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.961 0.505 1.303 0.595 ;
        RECT 0.225 0.735 1.051 0.825 ;
        RECT 0.961 0.505 1.051 0.825 ;
        RECT 0.25 0.735 0.355 0.975 ;
        RECT 0.225 0.685 0.34 0.825 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END S0
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.763 0.55 2.853 0.714 ;
        RECT 2.688 0.505 2.809 0.554 ;
        RECT 2.191 0.466 2.763 0.535 ;
        RECT 2.233 0.463 2.763 0.535 ;
        RECT 2.726 0.55 2.853 0.592 ;
        RECT 2.233 0.445 2.726 0.535 ;
        RECT 2.145 0.51 2.271 0.554 ;
        RECT 2.145 0.51 2.233 0.594 ;
        RECT 2.053 0.602 2.191 0.638 ;
        RECT 2.099 0.556 2.191 0.638 ;
        RECT 1.855 0.625 2.145 0.684 ;
        RECT 1.855 0.625 2.099 0.73 ;
        RECT 1.855 0.625 2.053 0.767 ;
        RECT 1.855 0.625 2.026 0.78 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.453 0.625 2.648 0.775 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.967 0.96 6.057 1.175 ;
      RECT 5.967 1.01 6.816 1.1 ;
      RECT 6.726 0.75 6.816 1.1 ;
      RECT 5.197 0.96 6.195 1.05 ;
      RECT 6.105 0.31 6.195 1.1 ;
      RECT 5.197 0.35 5.287 1.05 ;
      RECT 6.726 0.75 6.984 0.84 ;
      RECT 6.894 0.559 6.984 0.84 ;
      RECT 5.167 0.35 5.307 0.44 ;
      RECT 5.942 0.31 6.195 0.4 ;
      RECT 6.546 0.565 6.636 0.92 ;
      RECT 6.332 0.565 6.747 0.655 ;
      RECT 6.657 0.287 6.747 0.655 ;
      RECT 5.417 0.78 5.557 0.87 ;
      RECT 5.442 0.7 5.918 0.79 ;
      RECT 5.442 0.17 5.537 0.87 ;
      RECT 5.392 0.512 5.537 0.652 ;
      RECT 4.478 0.287 4.762 0.377 ;
      RECT 4.445 0.232 4.478 0.361 ;
      RECT 4.445 0.287 4.808 0.354 ;
      RECT 4.399 0.193 4.445 0.321 ;
      RECT 4.724 0.268 4.841 0.315 ;
      RECT 4.399 0.268 4.516 0.321 ;
      RECT 4.361 0.17 4.399 0.279 ;
      RECT 4.762 0.226 4.879 0.279 ;
      RECT 4.808 0.186 4.841 0.315 ;
      RECT 4.841 0.17 5.537 0.26 ;
      RECT 4.192 0.17 4.399 0.26 ;
      RECT 4.931 1.14 5.442 1.23 ;
      RECT 3.832 1.14 4.392 1.23 ;
      RECT 4.277 1.045 4.392 1.23 ;
      RECT 4.92 1.096 4.931 1.225 ;
      RECT 4.874 1.068 4.92 1.196 ;
      RECT 3.243 1.075 3.428 1.165 ;
      RECT 4.836 1.121 4.969 1.154 ;
      RECT 3.832 0.42 3.922 1.23 ;
      RECT 4.277 1.045 4.874 1.135 ;
      RECT 3.338 1.045 3.922 1.135 ;
      RECT 3.832 0.522 4.027 0.612 ;
      RECT 3.368 0.42 3.922 0.51 ;
      RECT 3.368 0.205 3.458 0.51 ;
      RECT 3.273 0.205 3.458 0.345 ;
      RECT 4.922 0.865 5.076 0.96 ;
      RECT 4.986 0.35 5.076 0.96 ;
      RECT 4.567 0.865 5.076 0.955 ;
      RECT 4.567 0.678 4.657 0.955 ;
      RECT 4.917 0.35 5.076 0.44 ;
      RECT 4.026 0.847 4.207 0.987 ;
      RECT 4.117 0.422 4.207 0.987 ;
      RECT 4.797 0.544 4.887 0.71 ;
      RECT 4.78 0.544 4.887 0.586 ;
      RECT 4.117 0.487 4.818 0.577 ;
      RECT 4.117 0.51 4.864 0.577 ;
      RECT 4.117 0.465 4.25 0.577 ;
      RECT 4.102 0.346 4.117 0.475 ;
      RECT 4.058 0.377 4.163 0.445 ;
      RECT 4.012 0.228 4.102 0.4 ;
      RECT 2.069 1.07 2.52 1.16 ;
      RECT 2.069 1.07 2.545 1.148 ;
      RECT 2.069 1.07 3.032 1.135 ;
      RECT 2.482 1.057 3.078 1.112 ;
      RECT 2.507 1.045 3.123 1.067 ;
      RECT 2.994 1.026 3.123 1.067 ;
      RECT 3.032 0.984 3.123 1.067 ;
      RECT 3.032 0.984 3.169 1.021 ;
      RECT 3.078 0.938 3.172 0.997 ;
      RECT 3.123 0.392 3.212 0.975 ;
      RECT 3.652 0.6 3.742 0.955 ;
      RECT 3.123 0.865 3.742 0.955 ;
      RECT 3.123 0.412 3.213 0.955 ;
      RECT 3.082 0.171 3.172 0.431 ;
      RECT 2.001 0.265 2.699 0.355 ;
      RECT 2.001 0.265 2.745 0.332 ;
      RECT 2.661 0.246 2.793 0.28 ;
      RECT 2.745 0.176 2.755 0.304 ;
      RECT 2.755 0.171 3.172 0.261 ;
      RECT 2.699 0.204 3.172 0.261 ;
      RECT 1.65 0.87 2.363 0.96 ;
      RECT 2.273 0.685 2.363 0.96 ;
      RECT 1.65 0.87 2.954 0.955 ;
      RECT 1.65 0.87 2.992 0.936 ;
      RECT 2.943 0.468 3.033 0.897 ;
      RECT 2.273 0.865 3.033 0.897 ;
      RECT 2.858 0.809 2.954 0.955 ;
      RECT 1.65 0.549 1.74 0.96 ;
      RECT 2.902 0.351 2.992 0.507 ;
      RECT 2.852 0.351 2.992 0.441 ;
      RECT 0.797 1.139 1.388 1.229 ;
      RECT 1.298 1.06 1.959 1.15 ;
      RECT 0.797 1.028 0.937 1.229 ;
      RECT 1.47 0.3 1.56 1.15 ;
      RECT 1.397 0.3 1.878 0.39 ;
      RECT 0.921 0.255 1.487 0.345 ;
      RECT 0.045 0.921 0.16 1.077 ;
      RECT 0.045 0.265 0.135 1.077 ;
      RECT 0.741 0.48 0.871 0.637 ;
      RECT 0.741 0.265 0.831 0.637 ;
      RECT 0.045 0.265 0.831 0.36 ;
  END
END MSDFFQX1H7R

MACRO MSDFFQX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MSDFFQX2H7R 0 0 ;
  SIZE 7.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7.6 1.48 ;
        RECT 7.397 0.834 7.537 1.48 ;
        RECT 6.906 0.93 6.996 1.48 ;
        RECT 6.441 1.23 6.581 1.48 ;
        RECT 5.707 1.225 5.852 1.48 ;
        RECT 4.657 1.225 4.797 1.48 ;
        RECT 3.508 1.225 3.648 1.48 ;
        RECT 2.593 1.225 2.733 1.48 ;
        RECT 1.478 1.24 1.618 1.48 ;
        RECT 0.304 1.092 0.444 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7.6 0.08 ;
        RECT 7.422 -0.08 7.512 0.466 ;
        RECT 6.922 -0.08 7.012 0.469 ;
        RECT 6.427 -0.08 6.517 0.425 ;
        RECT 5.712 -0.08 5.852 0.175 ;
        RECT 4.567 -0.08 4.707 0.175 ;
        RECT 3.548 -0.08 3.638 0.33 ;
        RECT 2.482 -0.08 2.622 0.175 ;
        RECT 1.563 -0.08 1.653 0.201 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.303 0.6 3.562 0.775 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END CK
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.455 0.609 0.645 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.189 0.71 1.38 0.97 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END D1
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.172 0.655 7.375 0.745 ;
        RECT 7.172 0.322 7.262 0.945 ;
      LAYER MET2 ;
        RECT 7.25 0.425 7.35 0.96 ;
      LAYER VIA1 ;
        RECT 7.255 0.655 7.345 0.745 ;
    END
  END Q
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.961 0.505 1.303 0.595 ;
        RECT 0.225 0.735 1.051 0.825 ;
        RECT 0.961 0.505 1.051 0.825 ;
        RECT 0.25 0.735 0.355 0.975 ;
        RECT 0.225 0.685 0.34 0.825 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END S0
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.763 0.55 2.853 0.714 ;
        RECT 2.688 0.505 2.809 0.554 ;
        RECT 2.191 0.466 2.763 0.535 ;
        RECT 2.233 0.463 2.763 0.535 ;
        RECT 2.726 0.55 2.853 0.592 ;
        RECT 2.233 0.445 2.726 0.535 ;
        RECT 2.145 0.51 2.271 0.554 ;
        RECT 2.145 0.51 2.233 0.594 ;
        RECT 2.053 0.602 2.191 0.638 ;
        RECT 2.099 0.556 2.191 0.638 ;
        RECT 1.855 0.625 2.145 0.684 ;
        RECT 1.855 0.625 2.099 0.73 ;
        RECT 1.855 0.625 2.053 0.767 ;
        RECT 1.855 0.625 2.026 0.78 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.453 0.685 2.673 0.775 ;
        RECT 2.453 0.625 2.638 0.775 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.967 0.96 6.057 1.175 ;
      RECT 5.967 1.01 6.816 1.1 ;
      RECT 6.726 0.75 6.816 1.1 ;
      RECT 5.197 0.96 6.195 1.05 ;
      RECT 6.105 0.31 6.195 1.1 ;
      RECT 5.197 0.35 5.287 1.05 ;
      RECT 6.726 0.75 6.984 0.84 ;
      RECT 6.894 0.559 6.984 0.84 ;
      RECT 5.167 0.35 5.307 0.44 ;
      RECT 5.942 0.31 6.195 0.4 ;
      RECT 6.546 0.565 6.636 0.92 ;
      RECT 6.332 0.565 6.747 0.655 ;
      RECT 6.657 0.287 6.747 0.655 ;
      RECT 5.417 0.78 5.557 0.87 ;
      RECT 5.442 0.7 5.918 0.79 ;
      RECT 5.442 0.17 5.537 0.87 ;
      RECT 5.392 0.512 5.537 0.652 ;
      RECT 4.456 0.265 4.784 0.355 ;
      RECT 4.445 0.221 4.456 0.35 ;
      RECT 4.445 0.265 4.83 0.332 ;
      RECT 4.399 0.193 4.445 0.321 ;
      RECT 4.746 0.246 4.879 0.279 ;
      RECT 4.83 0.175 4.841 0.304 ;
      RECT 4.361 0.246 4.494 0.279 ;
      RECT 4.841 0.17 5.537 0.26 ;
      RECT 4.192 0.17 4.399 0.26 ;
      RECT 4.784 0.204 5.537 0.26 ;
      RECT 4.931 1.14 5.442 1.23 ;
      RECT 3.832 1.14 4.392 1.23 ;
      RECT 4.277 1.045 4.392 1.23 ;
      RECT 4.92 1.096 4.931 1.225 ;
      RECT 4.874 1.068 4.92 1.196 ;
      RECT 3.243 1.075 3.428 1.165 ;
      RECT 4.836 1.121 4.969 1.154 ;
      RECT 3.832 0.42 3.922 1.23 ;
      RECT 4.277 1.045 4.874 1.135 ;
      RECT 3.338 1.045 3.922 1.135 ;
      RECT 3.832 0.522 4.027 0.612 ;
      RECT 3.368 0.42 3.922 0.51 ;
      RECT 3.368 0.205 3.458 0.51 ;
      RECT 3.273 0.205 3.458 0.345 ;
      RECT 4.922 0.865 5.076 0.96 ;
      RECT 4.986 0.35 5.076 0.96 ;
      RECT 4.567 0.865 5.076 0.955 ;
      RECT 4.567 0.678 4.657 0.955 ;
      RECT 4.917 0.35 5.076 0.44 ;
      RECT 4.026 0.847 4.207 0.987 ;
      RECT 4.117 0.422 4.207 0.987 ;
      RECT 4.797 0.545 4.887 0.71 ;
      RECT 4.782 0.545 4.887 0.587 ;
      RECT 4.117 0.489 4.82 0.579 ;
      RECT 4.117 0.512 4.866 0.579 ;
      RECT 4.117 0.466 4.252 0.579 ;
      RECT 4.102 0.346 4.117 0.475 ;
      RECT 4.058 0.377 4.163 0.445 ;
      RECT 4.012 0.228 4.102 0.4 ;
      RECT 2.069 1.07 2.52 1.16 ;
      RECT 2.069 1.07 2.545 1.148 ;
      RECT 2.069 1.07 3.032 1.135 ;
      RECT 2.482 1.057 3.078 1.112 ;
      RECT 2.507 1.045 3.123 1.067 ;
      RECT 2.994 1.026 3.123 1.067 ;
      RECT 3.032 0.984 3.123 1.067 ;
      RECT 3.032 0.984 3.169 1.021 ;
      RECT 3.078 0.938 3.172 0.997 ;
      RECT 3.123 0.392 3.212 0.975 ;
      RECT 3.652 0.6 3.742 0.955 ;
      RECT 3.123 0.865 3.742 0.955 ;
      RECT 3.123 0.412 3.213 0.955 ;
      RECT 3.082 0.171 3.172 0.431 ;
      RECT 2.001 0.265 2.699 0.355 ;
      RECT 2.001 0.265 2.745 0.332 ;
      RECT 2.661 0.246 2.793 0.28 ;
      RECT 2.745 0.176 2.755 0.304 ;
      RECT 2.755 0.171 3.172 0.261 ;
      RECT 2.699 0.204 3.172 0.261 ;
      RECT 1.65 0.87 2.363 0.96 ;
      RECT 2.273 0.685 2.363 0.96 ;
      RECT 1.65 0.87 2.954 0.955 ;
      RECT 1.65 0.87 2.992 0.936 ;
      RECT 2.943 0.468 3.033 0.897 ;
      RECT 2.273 0.865 3.033 0.897 ;
      RECT 2.858 0.809 2.954 0.955 ;
      RECT 1.65 0.549 1.74 0.96 ;
      RECT 2.902 0.351 2.992 0.507 ;
      RECT 2.852 0.351 2.992 0.441 ;
      RECT 0.847 1.139 1.388 1.229 ;
      RECT 1.298 1.06 1.959 1.15 ;
      RECT 0.847 1.028 0.937 1.229 ;
      RECT 0.797 1.028 0.937 1.118 ;
      RECT 1.47 0.3 1.56 1.15 ;
      RECT 1.397 0.3 1.56 0.41 ;
      RECT 1.397 0.3 1.878 0.39 ;
      RECT 0.921 0.255 1.487 0.345 ;
      RECT 0.045 0.921 0.16 1.077 ;
      RECT 0.045 0.265 0.135 1.077 ;
      RECT 0.741 0.48 0.871 0.637 ;
      RECT 0.741 0.265 0.831 0.637 ;
      RECT 0.045 0.265 0.831 0.36 ;
  END
END MSDFFQX2H7R

MACRO MSDFFQX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MSDFFQX3H7R 0 0 ;
  SIZE 7.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7.6 1.48 ;
        RECT 7.397 0.834 7.537 1.48 ;
        RECT 6.922 0.93 7.012 1.48 ;
        RECT 6.441 1.23 6.581 1.48 ;
        RECT 5.707 1.225 5.852 1.48 ;
        RECT 4.657 1.225 4.797 1.48 ;
        RECT 3.508 1.225 3.648 1.48 ;
        RECT 2.593 1.225 2.733 1.48 ;
        RECT 1.478 1.24 1.618 1.48 ;
        RECT 0.304 1.092 0.444 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7.6 0.08 ;
        RECT 7.422 -0.08 7.512 0.466 ;
        RECT 6.922 -0.08 7.012 0.391 ;
        RECT 6.427 -0.08 6.517 0.425 ;
        RECT 5.712 -0.08 5.852 0.175 ;
        RECT 4.567 -0.08 4.707 0.175 ;
        RECT 3.548 -0.08 3.638 0.33 ;
        RECT 2.482 -0.08 2.622 0.175 ;
        RECT 1.563 -0.08 1.653 0.201 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.303 0.6 3.562 0.775 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END CK
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.455 0.609 0.645 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.178 0.844 1.379 0.97 ;
        RECT 1.221 0.71 1.379 0.97 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END D1
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.172 0.655 7.375 0.745 ;
        RECT 7.172 0.322 7.262 0.945 ;
      LAYER MET2 ;
        RECT 7.25 0.425 7.35 0.96 ;
      LAYER VIA1 ;
        RECT 7.255 0.655 7.345 0.745 ;
    END
  END Q
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.961 0.505 1.303 0.595 ;
        RECT 0.225 0.735 1.051 0.825 ;
        RECT 0.961 0.505 1.051 0.825 ;
        RECT 0.25 0.735 0.355 0.98 ;
        RECT 0.225 0.685 0.34 0.825 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END S0
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.763 0.55 2.853 0.714 ;
        RECT 2.688 0.505 2.809 0.554 ;
        RECT 2.191 0.466 2.763 0.535 ;
        RECT 2.233 0.463 2.763 0.535 ;
        RECT 2.726 0.55 2.853 0.592 ;
        RECT 2.233 0.445 2.726 0.535 ;
        RECT 2.145 0.51 2.271 0.554 ;
        RECT 2.145 0.51 2.233 0.594 ;
        RECT 2.053 0.602 2.191 0.638 ;
        RECT 2.099 0.556 2.191 0.638 ;
        RECT 1.855 0.625 2.145 0.684 ;
        RECT 1.855 0.625 2.099 0.73 ;
        RECT 1.855 0.625 2.053 0.767 ;
        RECT 1.855 0.625 2.026 0.78 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.453 0.625 2.648 0.775 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.967 0.96 6.057 1.175 ;
      RECT 5.967 1.01 6.832 1.1 ;
      RECT 6.742 0.75 6.832 1.1 ;
      RECT 5.197 0.96 6.195 1.05 ;
      RECT 6.105 0.31 6.195 1.1 ;
      RECT 5.197 0.35 5.287 1.05 ;
      RECT 6.742 0.75 6.984 0.84 ;
      RECT 6.894 0.559 6.984 0.84 ;
      RECT 5.167 0.35 5.307 0.44 ;
      RECT 5.942 0.31 6.195 0.4 ;
      RECT 6.546 0.565 6.636 0.92 ;
      RECT 6.332 0.565 6.747 0.655 ;
      RECT 6.657 0.287 6.747 0.655 ;
      RECT 5.417 0.78 5.557 0.87 ;
      RECT 5.442 0.7 5.918 0.79 ;
      RECT 5.442 0.17 5.532 0.87 ;
      RECT 5.392 0.512 5.532 0.652 ;
      RECT 5.442 0.17 5.537 0.425 ;
      RECT 4.509 0.318 4.731 0.408 ;
      RECT 4.491 0.271 4.509 0.399 ;
      RECT 4.491 0.318 4.777 0.385 ;
      RECT 4.445 0.239 4.491 0.367 ;
      RECT 4.399 0.193 4.445 0.321 ;
      RECT 4.693 0.299 4.823 0.339 ;
      RECT 4.399 0.299 4.547 0.321 ;
      RECT 4.731 0.257 4.841 0.307 ;
      RECT 4.731 0.257 4.879 0.279 ;
      RECT 4.361 0.17 4.399 0.279 ;
      RECT 4.841 0.17 5.537 0.26 ;
      RECT 4.192 0.17 4.399 0.26 ;
      RECT 4.777 0.211 5.537 0.26 ;
      RECT 4.823 0.179 4.841 0.307 ;
      RECT 4.931 1.14 5.442 1.23 ;
      RECT 3.832 1.14 4.392 1.23 ;
      RECT 4.277 1.045 4.392 1.23 ;
      RECT 4.92 1.096 4.931 1.225 ;
      RECT 4.874 1.068 4.92 1.196 ;
      RECT 3.243 1.075 3.428 1.165 ;
      RECT 4.836 1.121 4.969 1.154 ;
      RECT 3.832 0.42 3.922 1.23 ;
      RECT 4.277 1.045 4.874 1.135 ;
      RECT 3.338 1.045 3.922 1.135 ;
      RECT 3.832 0.522 4.027 0.612 ;
      RECT 3.368 0.42 3.922 0.51 ;
      RECT 3.368 0.205 3.458 0.51 ;
      RECT 3.273 0.205 3.458 0.345 ;
      RECT 4.922 0.865 5.076 0.96 ;
      RECT 4.986 0.35 5.076 0.96 ;
      RECT 4.567 0.865 5.076 0.955 ;
      RECT 4.567 0.678 4.657 0.955 ;
      RECT 4.917 0.35 5.076 0.44 ;
      RECT 4.026 0.847 4.207 0.987 ;
      RECT 4.117 0.422 4.207 0.987 ;
      RECT 4.797 0.55 4.887 0.71 ;
      RECT 4.791 0.55 4.887 0.591 ;
      RECT 4.117 0.498 4.829 0.588 ;
      RECT 4.117 0.521 4.875 0.588 ;
      RECT 4.117 0.494 4.261 0.588 ;
      RECT 4.117 0.467 4.253 0.588 ;
      RECT 4.102 0.346 4.117 0.475 ;
      RECT 4.058 0.377 4.163 0.445 ;
      RECT 4.012 0.228 4.102 0.4 ;
      RECT 2.069 1.08 2.51 1.17 ;
      RECT 2.069 1.08 2.545 1.153 ;
      RECT 2.069 1.08 3.032 1.135 ;
      RECT 2.472 1.062 3.078 1.112 ;
      RECT 2.507 1.045 3.123 1.067 ;
      RECT 2.994 1.026 3.123 1.067 ;
      RECT 3.032 0.984 3.123 1.067 ;
      RECT 3.032 0.984 3.169 1.021 ;
      RECT 3.078 0.938 3.172 0.997 ;
      RECT 3.123 0.392 3.212 0.975 ;
      RECT 3.652 0.6 3.742 0.955 ;
      RECT 3.123 0.865 3.742 0.955 ;
      RECT 3.123 0.412 3.213 0.955 ;
      RECT 3.082 0.171 3.172 0.431 ;
      RECT 2.001 0.265 2.699 0.355 ;
      RECT 2.001 0.265 2.745 0.332 ;
      RECT 2.661 0.246 2.793 0.28 ;
      RECT 2.745 0.176 2.755 0.304 ;
      RECT 2.755 0.171 3.172 0.261 ;
      RECT 2.699 0.204 3.172 0.261 ;
      RECT 1.65 0.87 2.363 0.96 ;
      RECT 2.273 0.685 2.363 0.96 ;
      RECT 1.65 0.87 2.954 0.955 ;
      RECT 1.65 0.87 2.992 0.936 ;
      RECT 2.943 0.468 3.033 0.897 ;
      RECT 2.273 0.865 3.033 0.897 ;
      RECT 2.858 0.809 2.954 0.955 ;
      RECT 1.65 0.549 1.74 0.96 ;
      RECT 2.902 0.351 2.992 0.507 ;
      RECT 2.852 0.351 2.992 0.441 ;
      RECT 0.847 1.139 1.388 1.229 ;
      RECT 1.298 1.06 1.959 1.15 ;
      RECT 0.847 1.028 0.937 1.229 ;
      RECT 0.797 1.028 0.937 1.118 ;
      RECT 1.47 0.3 1.56 1.15 ;
      RECT 1.397 0.3 1.56 0.41 ;
      RECT 1.397 0.3 1.878 0.39 ;
      RECT 0.921 0.252 1.487 0.342 ;
      RECT 0.045 0.921 0.16 1.061 ;
      RECT 0.045 0.265 0.135 1.061 ;
      RECT 0.741 0.48 0.871 0.637 ;
      RECT 0.741 0.265 0.831 0.637 ;
      RECT 0.045 0.265 0.831 0.355 ;
  END
END MSDFFQX3H7R

MACRO MUX2X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2X0P5H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.49 0.95 1.58 1.48 ;
        RECT 0.31 1.045 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.56 -0.08 1.65 0.33 ;
        RECT 0.295 -0.08 0.435 0.325 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.595 0.6 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.41 0.425 1.635 0.545 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END B
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.23 0.17 1.32 0.555 ;
        RECT 0.66 0.17 1.32 0.26 ;
        RECT 0.25 0.415 0.75 0.505 ;
        RECT 0.66 0.17 0.75 0.505 ;
        RECT 0.25 0.415 0.345 0.58 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.715 0.935 1.945 1.025 ;
        RECT 1.855 0.23 1.945 1.025 ;
        RECT 1.785 0.23 1.945 0.32 ;
      LAYER MET2 ;
        RECT 1.85 0.225 1.95 0.76 ;
      LAYER VIA1 ;
        RECT 1.855 0.455 1.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.81 0.725 0.9 0.94 ;
      RECT 0.81 0.725 1.755 0.815 ;
      RECT 1.045 0.35 1.135 0.815 ;
      RECT 0.995 0.35 1.135 0.44 ;
      RECT 0.54 1.09 1.025 1.18 ;
      RECT 0.54 0.865 0.63 1.18 ;
      RECT 0.07 0.865 0.63 0.955 ;
      RECT 0.07 0.225 0.16 0.955 ;
  END
END MUX2X0P5H7R

MACRO MUX2X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2X0P7H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.49 0.982 1.58 1.48 ;
        RECT 0.31 1.045 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.56 -0.08 1.65 0.33 ;
        RECT 0.295 -0.08 0.435 0.325 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.595 0.6 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.41 0.425 1.635 0.545 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END B
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.23 0.17 1.32 0.555 ;
        RECT 0.66 0.17 1.32 0.26 ;
        RECT 0.25 0.415 0.75 0.505 ;
        RECT 0.66 0.17 0.75 0.505 ;
        RECT 0.25 0.415 0.345 0.58 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.715 0.935 1.945 1.025 ;
        RECT 1.855 0.254 1.945 1.025 ;
        RECT 1.785 0.254 1.945 0.344 ;
      LAYER MET2 ;
        RECT 1.85 0.225 1.95 0.76 ;
      LAYER VIA1 ;
        RECT 1.855 0.455 1.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.81 0.725 0.9 0.94 ;
      RECT 0.81 0.725 1.755 0.815 ;
      RECT 1.045 0.35 1.135 0.815 ;
      RECT 0.995 0.35 1.135 0.44 ;
      RECT 0.54 1.09 1.025 1.18 ;
      RECT 0.54 0.865 0.63 1.18 ;
      RECT 0.07 0.865 0.63 0.955 ;
      RECT 0.07 0.21 0.16 0.955 ;
  END
END MUX2X0P7H7R

MACRO MUX2X12H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2X12H7R 0 0 ;
  SIZE 6.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.4 1.48 ;
        RECT 5.826 1.05 5.916 1.48 ;
        RECT 5.326 1.05 5.416 1.48 ;
        RECT 4.826 1.05 4.916 1.48 ;
        RECT 4.274 1.225 4.414 1.48 ;
        RECT 3.714 1.24 3.854 1.48 ;
        RECT 1.107 1.24 1.247 1.48 ;
        RECT 0.585 1.05 0.675 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.4 0.08 ;
        RECT 5.674 -0.08 5.814 0.307 ;
        RECT 5.174 -0.08 5.314 0.307 ;
        RECT 4.674 -0.08 4.814 0.306 ;
        RECT 4.026 -0.08 4.166 0.161 ;
        RECT 3.332 -0.08 3.472 0.161 ;
        RECT 1.107 -0.08 1.247 0.205 ;
        RECT 0.585 -0.08 0.675 0.35 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.76 0.655 1.3 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.584 0.655 3.924 0.745 ;
      LAYER MET2 ;
        RECT 3.65 0.43 3.75 0.96 ;
      LAYER VIA1 ;
        RECT 3.655 0.655 3.745 0.745 ;
    END
  END B
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.39 0.735 1.889 0.825 ;
        RECT 0.475 0.855 1.48 0.945 ;
        RECT 1.39 0.735 1.48 0.945 ;
        RECT 0.475 0.726 0.565 0.945 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.076 0.866 6.166 1.006 ;
        RECT 4.576 0.866 6.166 0.956 ;
        RECT 4.449 0.402 6.039 0.492 ;
        RECT 5.949 0.31 6.039 0.492 ;
        RECT 5.855 0.402 5.945 0.956 ;
        RECT 5.576 0.866 5.666 1.006 ;
        RECT 5.449 0.325 5.539 0.492 ;
        RECT 5.076 0.866 5.166 1.006 ;
        RECT 4.949 0.325 5.039 0.492 ;
        RECT 4.576 0.866 4.666 1.006 ;
        RECT 4.449 0.336 4.539 0.492 ;
      LAYER MET2 ;
        RECT 5.85 0.43 5.95 0.96 ;
      LAYER VIA1 ;
        RECT 5.855 0.655 5.945 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.742 1.14 3.558 1.23 ;
      RECT 3.676 1.06 4.18 1.15 ;
      RECT 4.396 0.656 5.621 0.746 ;
      RECT 3.292 0.251 3.512 0.341 ;
      RECT 1.667 0.171 3.174 0.261 ;
      RECT 3.631 0.17 3.867 0.26 ;
      RECT 4.391 0.656 4.396 0.975 ;
      RECT 4.352 0.636 4.391 0.997 ;
      RECT 4.306 0.594 4.352 1.039 ;
      RECT 4.273 0.554 4.306 0.683 ;
      RECT 4.227 0.515 4.273 0.643 ;
      RECT 4.181 0.469 4.227 0.597 ;
      RECT 4.135 0.423 4.181 0.551 ;
      RECT 4.089 0.377 4.135 0.505 ;
      RECT 4.043 0.331 4.089 0.459 ;
      RECT 3.997 0.285 4.043 0.413 ;
      RECT 3.951 0.239 3.997 0.367 ;
      RECT 3.905 0.193 3.951 0.321 ;
      RECT 4.264 0.955 4.306 1.083 ;
      RECT 4.218 0.999 4.264 1.127 ;
      RECT 4.18 1.041 4.218 1.15 ;
      RECT 3.867 0.17 3.905 0.279 ;
      RECT 3.638 1.06 3.676 1.169 ;
      RECT 3.596 1.081 3.638 1.209 ;
      RECT 3.593 0.17 3.631 0.279 ;
      RECT 3.558 1.121 3.596 1.23 ;
      RECT 3.55 0.191 3.593 0.32 ;
      RECT 3.512 0.232 3.55 0.341 ;
      RECT 3.254 0.232 3.292 0.341 ;
      RECT 3.212 0.192 3.254 0.32 ;
      RECT 3.174 0.171 3.212 0.28 ;
      RECT 2.874 0.95 3.519 1.04 ;
      RECT 3.429 0.88 4.134 0.97 ;
      RECT 3.044 0.351 3.134 1.04 ;
      RECT 3.044 0.431 3.834 0.521 ;
      RECT 3.694 0.356 3.834 0.521 ;
      RECT 2.462 0.351 3.134 0.441 ;
      RECT 0.827 1.06 1.558 1.15 ;
      RECT 0.827 1.06 1.604 1.127 ;
      RECT 0.827 1.06 1.62 1.096 ;
      RECT 1.52 1.041 1.658 1.069 ;
      RECT 1.558 0.999 2.65 1.05 ;
      RECT 1.604 0.968 2.702 1.001 ;
      RECT 2.702 0.531 2.748 0.975 ;
      RECT 1.62 0.96 2.748 0.975 ;
      RECT 2.696 0.873 2.702 1.001 ;
      RECT 2.612 0.941 2.748 0.975 ;
      RECT 2.65 0.899 2.696 1.027 ;
      RECT 2.702 0.531 2.792 0.93 ;
      RECT 2.224 0.531 2.792 0.621 ;
      RECT 2.22 0.491 2.224 0.619 ;
      RECT 2.174 0.466 2.22 0.594 ;
      RECT 2.128 0.42 2.174 0.548 ;
      RECT 2.128 0.512 2.262 0.548 ;
      RECT 2.082 0.374 2.128 0.502 ;
      RECT 2.044 0.42 2.174 0.46 ;
      RECT 1.589 0.351 2.082 0.441 ;
      RECT 1.571 0.304 1.589 0.432 ;
      RECT 1.533 0.374 2.128 0.404 ;
      RECT 0.827 0.295 1.571 0.385 ;
      RECT 0.827 0.332 1.627 0.385 ;
      RECT 0.295 1.026 0.435 1.116 ;
      RECT 0.295 0.256 0.385 1.116 ;
      RECT 2.125 0.74 2.612 0.83 ;
      RECT 2.097 0.688 2.125 0.816 ;
      RECT 2.051 0.651 2.097 0.779 ;
      RECT 2.051 0.721 2.163 0.779 ;
      RECT 2.005 0.605 2.051 0.733 ;
      RECT 1.959 0.559 2.005 0.687 ;
      RECT 1.921 0.605 2.051 0.645 ;
      RECT 1.487 0.536 1.959 0.626 ;
      RECT 1.464 0.486 1.487 0.615 ;
      RECT 1.426 0.559 2.005 0.584 ;
      RECT 0.295 0.475 1.464 0.565 ;
      RECT 0.295 0.517 1.525 0.565 ;
      RECT 0.295 0.256 0.435 0.346 ;
  END
END MUX2X12H7R

MACRO MUX2X16H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2X16H7R 0 0 ;
  SIZE 9 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 9 1.48 ;
        RECT 8.833 1.035 8.923 1.48 ;
        RECT 8.308 1.075 8.448 1.48 ;
        RECT 7.778 1.061 7.918 1.48 ;
        RECT 7.263 1.075 7.403 1.48 ;
        RECT 6.763 1.075 6.903 1.48 ;
        RECT 6.273 1.2 6.363 1.48 ;
        RECT 5.71 1.24 5.85 1.48 ;
        RECT 5.15 1.24 5.29 1.48 ;
        RECT 1.632 1.215 1.772 1.48 ;
        RECT 1.072 1.215 1.212 1.48 ;
        RECT 0.585 1.035 0.675 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 9 0.08 ;
        RECT 8.724 -0.08 8.814 0.36 ;
        RECT 8.199 -0.08 8.339 0.32 ;
        RECT 7.699 -0.08 7.839 0.32 ;
        RECT 7.199 -0.08 7.339 0.32 ;
        RECT 6.699 -0.08 6.839 0.32 ;
        RECT 6.169 -0.08 6.309 0.16 ;
        RECT 5.494 -0.08 5.634 0.16 ;
        RECT 4.768 -0.08 4.908 0.16 ;
        RECT 1.632 -0.08 1.772 0.205 ;
        RECT 1.072 -0.08 1.212 0.205 ;
        RECT 0.585 -0.08 0.675 0.365 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.972 0.655 1.712 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.978 0.65 5.918 0.745 ;
      LAYER MET2 ;
        RECT 5.25 0.425 5.35 0.96 ;
      LAYER VIA1 ;
        RECT 5.255 0.655 5.345 0.745 ;
    END
  END B
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.986 0.777 2.763 0.867 ;
        RECT 0.5 0.855 2.024 0.886 ;
        RECT 1.908 0.836 2.763 0.867 ;
        RECT 1.946 0.797 1.986 0.925 ;
        RECT 0.5 0.855 1.946 0.945 ;
        RECT 0.5 0.805 0.59 0.945 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 8.583 0.881 8.673 1.021 ;
        RECT 6.538 0.881 8.673 0.971 ;
        RECT 6.474 0.41 8.564 0.5 ;
        RECT 8.474 0.325 8.564 0.5 ;
        RECT 8.455 0.41 8.545 0.971 ;
        RECT 8.068 0.881 8.158 1.021 ;
        RECT 7.974 0.325 8.064 0.5 ;
        RECT 7.538 0.881 7.628 1.021 ;
        RECT 7.474 0.325 7.564 0.5 ;
        RECT 7.038 0.881 7.128 1.021 ;
        RECT 6.974 0.325 7.064 0.5 ;
        RECT 6.538 0.881 6.628 1.021 ;
        RECT 6.474 0.325 6.564 0.5 ;
      LAYER MET2 ;
        RECT 8.45 0.43 8.55 0.96 ;
      LAYER VIA1 ;
        RECT 8.455 0.655 8.545 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.19 1.14 4.993 1.23 ;
      RECT 5.111 1.06 6.15 1.15 ;
      RECT 6.384 0.59 8.365 0.68 ;
      RECT 4.635 0.251 4.975 0.341 ;
      RECT 5.455 0.25 5.672 0.34 ;
      RECT 5.775 0.185 6.028 0.275 ;
      RECT 5.079 0.185 5.352 0.275 ;
      RECT 2.19 0.17 4.516 0.26 ;
      RECT 6.34 0.481 6.384 0.976 ;
      RECT 6.294 0.436 6.34 1.021 ;
      RECT 6.25 0.391 6.294 0.519 ;
      RECT 6.204 0.346 6.25 0.474 ;
      RECT 6.158 0.3 6.204 0.428 ;
      RECT 6.112 0.254 6.158 0.382 ;
      RECT 6.066 0.208 6.112 0.336 ;
      RECT 6.28 0.923 6.294 1.051 ;
      RECT 6.234 0.953 6.28 1.081 ;
      RECT 6.188 0.999 6.234 1.127 ;
      RECT 6.15 1.041 6.188 1.15 ;
      RECT 6.028 0.185 6.066 0.294 ;
      RECT 5.737 0.185 5.775 0.294 ;
      RECT 5.71 0.198 5.737 0.327 ;
      RECT 5.672 0.231 5.71 0.34 ;
      RECT 5.417 0.231 5.455 0.34 ;
      RECT 5.39 0.198 5.417 0.327 ;
      RECT 5.352 0.185 5.39 0.294 ;
      RECT 5.073 1.06 5.111 1.169 ;
      RECT 5.041 0.185 5.079 0.294 ;
      RECT 5.031 1.081 5.073 1.209 ;
      RECT 5.013 0.199 5.041 0.327 ;
      RECT 4.993 1.121 5.031 1.23 ;
      RECT 4.975 0.232 5.013 0.341 ;
      RECT 4.597 0.232 4.635 0.341 ;
      RECT 4.554 0.191 4.597 0.32 ;
      RECT 4.516 0.17 4.554 0.279 ;
      RECT 3.755 0.947 4.955 1.037 ;
      RECT 3.755 0.947 6.073 0.97 ;
      RECT 4.865 0.88 6.118 0.948 ;
      RECT 3.755 0.35 3.845 1.037 ;
      RECT 6.03 0.785 6.12 0.925 ;
      RECT 4.388 0.431 5.97 0.521 ;
      RECT 5.83 0.365 5.97 0.521 ;
      RECT 3.253 0.35 4.478 0.44 ;
      RECT 5.157 0.365 5.297 0.521 ;
      RECT 0.787 1.035 2.077 1.125 ;
      RECT 0.787 1.035 2.115 1.106 ;
      RECT 0.787 1.035 2.152 1.069 ;
      RECT 0.787 1.035 3.551 1.05 ;
      RECT 2.039 1.016 3.575 1.038 ;
      RECT 2.077 0.978 3.575 1.038 ;
      RECT 2.115 0.96 3.621 1.003 ;
      RECT 3.551 0.91 3.575 1.038 ;
      RECT 3.513 0.941 3.621 1.003 ;
      RECT 2.115 0.959 2.154 1.05 ;
      RECT 3.575 0.53 3.665 0.958 ;
      RECT 3.048 0.53 3.665 0.62 ;
      RECT 3.048 0.35 3.138 0.62 ;
      RECT 2.113 0.35 3.138 0.44 ;
      RECT 2.096 0.303 2.113 0.432 ;
      RECT 2.058 0.35 3.138 0.404 ;
      RECT 0.792 0.295 2.096 0.385 ;
      RECT 0.792 0.331 2.151 0.385 ;
      RECT 0.32 0.24 0.41 1.12 ;
      RECT 2.858 0.77 3.485 0.86 ;
      RECT 2.858 0.546 2.948 0.86 ;
      RECT 1.963 0.546 2.948 0.636 ;
      RECT 1.93 0.491 1.963 0.62 ;
      RECT 1.892 0.546 2.948 0.584 ;
      RECT 0.32 0.475 1.93 0.565 ;
      RECT 0.32 0.527 2.001 0.565 ;
  END
END MUX2X16H7R

MACRO MUX2X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2X1H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.49 1.03 1.58 1.48 ;
        RECT 0.31 1.045 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.56 -0.08 1.65 0.33 ;
        RECT 0.295 -0.08 0.435 0.325 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.595 0.6 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.41 0.425 1.635 0.545 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END B
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.23 0.17 1.32 0.555 ;
        RECT 0.66 0.17 1.32 0.26 ;
        RECT 0.25 0.415 0.75 0.505 ;
        RECT 0.66 0.17 0.75 0.505 ;
        RECT 0.25 0.415 0.345 0.58 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.715 0.935 1.945 1.025 ;
        RECT 1.855 0.29 1.945 1.025 ;
        RECT 1.785 0.29 1.945 0.38 ;
      LAYER MET2 ;
        RECT 1.85 0.225 1.95 0.76 ;
      LAYER VIA1 ;
        RECT 1.855 0.455 1.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.81 0.725 0.9 0.94 ;
      RECT 0.81 0.725 1.755 0.815 ;
      RECT 1.045 0.35 1.135 0.815 ;
      RECT 0.995 0.35 1.135 0.44 ;
      RECT 0.54 1.09 1.025 1.18 ;
      RECT 0.54 0.865 0.63 1.18 ;
      RECT 0.07 0.865 0.63 0.955 ;
      RECT 0.07 0.225 0.16 0.955 ;
  END
END MUX2X1H7R

MACRO MUX2X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2X1P4H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.49 1.055 1.58 1.48 ;
        RECT 0.31 1.045 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.56 -0.08 1.65 0.33 ;
        RECT 0.295 -0.08 0.435 0.325 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.595 0.6 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.41 0.425 1.635 0.545 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END B
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.23 0.17 1.32 0.555 ;
        RECT 0.66 0.17 1.32 0.26 ;
        RECT 0.25 0.415 0.75 0.505 ;
        RECT 0.66 0.17 0.75 0.505 ;
        RECT 0.25 0.415 0.345 0.58 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.715 0.916 1.945 1.006 ;
        RECT 1.855 0.326 1.945 1.006 ;
        RECT 1.785 0.326 1.945 0.416 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.81 0.706 0.9 0.94 ;
      RECT 0.81 0.706 1.757 0.796 ;
      RECT 1.045 0.35 1.135 0.796 ;
      RECT 0.995 0.35 1.135 0.44 ;
      RECT 0.54 1.09 1.025 1.18 ;
      RECT 0.54 0.865 0.63 1.18 ;
      RECT 0.07 0.865 0.63 0.955 ;
      RECT 0.07 0.22 0.16 0.955 ;
  END
END MUX2X1P4H7R

MACRO MUX2X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2X2H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 2.29 1.035 2.38 1.48 ;
        RECT 1.775 1.165 1.865 1.48 ;
        RECT 0.31 1.225 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 2.29 -0.08 2.38 0.365 ;
        RECT 1.73 -0.08 1.82 0.35 ;
        RECT 0.31 -0.08 0.45 0.325 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.405 0.595 0.585 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.58 0.625 1.78 0.76 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.685 0.725 0.775 0.884 ;
        RECT 0.225 0.855 0.745 0.922 ;
        RECT 0.225 0.855 0.699 0.945 ;
        RECT 0.661 0.843 0.775 0.884 ;
        RECT 0.225 0.785 0.315 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.015 1.075 2.18 1.165 ;
        RECT 2.09 0.255 2.18 1.165 ;
        RECT 2.015 0.255 2.18 0.345 ;
      LAYER MET2 ;
        RECT 2.05 0.18 2.15 0.56 ;
      LAYER VIA1 ;
        RECT 2.055 0.255 2.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.23 1.04 1.32 1.18 ;
      RECT 1.23 1.04 1.678 1.13 ;
      RECT 1.23 1.04 1.724 1.107 ;
      RECT 1.64 1.021 1.77 1.061 ;
      RECT 1.678 0.979 1.77 1.061 ;
      RECT 1.724 0.933 1.816 1.015 ;
      RECT 1.77 0.887 1.862 0.969 ;
      RECT 1.77 0.887 1.908 0.923 ;
      RECT 1.816 0.841 1.91 0.899 ;
      RECT 1.862 0.795 1.956 0.875 ;
      RECT 1.908 0.771 1.91 0.899 ;
      RECT 1.91 0.44 2 0.83 ;
      RECT 1.535 0.44 2 0.53 ;
      RECT 1.535 0.17 1.625 0.53 ;
      RECT 1.05 0.17 1.14 0.35 ;
      RECT 1.05 0.17 1.625 0.26 ;
      RECT 1.4 0.85 1.61 0.94 ;
      RECT 1.4 0.63 1.49 0.94 ;
      RECT 1.305 0.63 1.49 0.72 ;
      RECT 1.305 0.35 1.395 0.72 ;
      RECT 1.305 0.35 1.445 0.44 ;
      RECT 0.54 1.14 1.14 1.23 ;
      RECT 1.05 0.86 1.14 1.23 ;
      RECT 0.54 1.04 0.63 1.23 ;
      RECT 0.045 1.04 0.63 1.13 ;
      RECT 0.045 0.225 0.135 1.13 ;
      RECT 1.05 0.86 1.31 0.95 ;
      RECT 1.22 0.81 1.31 0.95 ;
      RECT 0.69 0.415 0.78 0.575 ;
      RECT 0.045 0.415 0.78 0.505 ;
      RECT 0.045 0.225 0.16 0.505 ;
      RECT 0.82 0.96 0.96 1.05 ;
      RECT 0.87 0.235 0.96 1.05 ;
      RECT 0.575 0.235 0.96 0.325 ;
  END
END MUX2X2H7R

MACRO MUX2X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2X3H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 2.292 1.035 2.382 1.48 ;
        RECT 1.752 1.225 1.892 1.48 ;
        RECT 0.31 1.225 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 2.293 -0.08 2.383 0.365 ;
        RECT 1.792 -0.08 1.882 0.35 ;
        RECT 0.31 -0.08 0.45 0.325 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.415 0.615 0.595 0.765 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.605 0.62 1.755 0.8 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.855 0.78 0.945 ;
        RECT 0.69 0.739 0.78 0.945 ;
        RECT 0.225 0.775 0.315 0.945 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.017 0.96 2.175 1.05 ;
        RECT 2.085 0.255 2.175 1.05 ;
        RECT 2.017 0.255 2.175 0.345 ;
      LAYER MET2 ;
        RECT 2.05 0.18 2.15 0.56 ;
      LAYER VIA1 ;
        RECT 2.055 0.255 2.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.23 1.1 1.658 1.19 ;
      RECT 1.23 1.1 1.704 1.167 ;
      RECT 1.62 1.081 1.75 1.121 ;
      RECT 1.23 1.05 1.321 1.19 ;
      RECT 1.658 1.039 1.75 1.121 ;
      RECT 1.704 0.993 1.796 1.075 ;
      RECT 1.75 0.947 1.842 1.029 ;
      RECT 1.75 0.947 1.888 0.983 ;
      RECT 1.796 0.901 1.905 0.952 ;
      RECT 1.842 0.855 1.951 0.92 ;
      RECT 1.888 0.823 1.905 0.952 ;
      RECT 1.905 0.44 1.995 0.875 ;
      RECT 1.605 0.44 1.995 0.53 ;
      RECT 1.605 0.17 1.702 0.53 ;
      RECT 1.08 0.17 1.17 0.36 ;
      RECT 1.08 0.17 1.702 0.26 ;
      RECT 1.425 0.89 1.61 0.98 ;
      RECT 1.425 0.35 1.515 0.98 ;
      RECT 1.335 0.35 1.515 0.44 ;
      RECT 0.54 1.14 1.14 1.23 ;
      RECT 1.05 0.81 1.14 1.23 ;
      RECT 0.54 1.04 0.63 1.23 ;
      RECT 0.045 1.04 0.63 1.13 ;
      RECT 0.045 0.235 0.135 1.13 ;
      RECT 1.05 0.81 1.335 0.9 ;
      RECT 1.245 0.75 1.335 0.9 ;
      RECT 0.72 0.435 0.81 0.6 ;
      RECT 0.045 0.435 0.81 0.525 ;
      RECT 0.045 0.235 0.16 0.525 ;
      RECT 0.87 0.696 0.96 1.05 ;
      RECT 0.9 0.255 0.99 0.734 ;
      RECT 0.645 0.255 0.99 0.345 ;
  END
END MUX2X3H7R

MACRO MUX2X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2X4H7R 0 0 ;
  SIZE 2.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.8 1.48 ;
        RECT 2.325 1.05 2.415 1.48 ;
        RECT 1.785 1.225 1.925 1.48 ;
        RECT 0.31 1.215 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.8 0.08 ;
        RECT 2.32 -0.08 2.41 0.35 ;
        RECT 1.82 -0.08 1.91 0.35 ;
        RECT 0.335 -0.08 0.425 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.405 0.63 0.605 0.765 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.64 0.625 1.82 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.855 0.795 0.945 ;
        RECT 0.705 0.738 0.795 0.945 ;
        RECT 0.225 0.765 0.315 0.945 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.575 0.275 2.665 1.075 ;
        RECT 2.105 0.655 2.665 0.745 ;
        RECT 2.05 0.965 2.195 1.055 ;
        RECT 2.105 0.26 2.195 1.055 ;
        RECT 2.045 0.26 2.195 0.35 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.265 1.055 1.738 1.145 ;
      RECT 1.265 1.055 1.784 1.122 ;
      RECT 1.7 1.036 1.83 1.076 ;
      RECT 1.265 1.005 1.356 1.145 ;
      RECT 1.738 0.994 1.83 1.076 ;
      RECT 1.784 0.948 1.876 1.03 ;
      RECT 1.83 0.902 1.92 0.985 ;
      RECT 1.876 0.857 1.966 0.94 ;
      RECT 1.92 0.44 2.01 0.895 ;
      RECT 1.64 0.44 2.01 0.53 ;
      RECT 1.64 0.17 1.73 0.53 ;
      RECT 1.085 0.17 1.175 0.33 ;
      RECT 1.085 0.17 1.73 0.26 ;
      RECT 1.46 0.875 1.66 0.965 ;
      RECT 1.46 0.35 1.55 0.965 ;
      RECT 1.375 0.35 1.55 0.44 ;
      RECT 0.54 1.14 1.175 1.23 ;
      RECT 1.085 0.81 1.175 1.23 ;
      RECT 0.54 1.035 0.63 1.23 ;
      RECT 0.045 1.035 0.63 1.125 ;
      RECT 0.045 0.25 0.135 1.125 ;
      RECT 1.085 0.81 1.37 0.9 ;
      RECT 1.28 0.71 1.37 0.9 ;
      RECT 0.72 0.45 0.81 0.63 ;
      RECT 0.045 0.45 0.81 0.54 ;
      RECT 0.045 0.25 0.185 0.34 ;
      RECT 0.905 0.27 0.995 1.035 ;
      RECT 0.625 0.27 0.995 0.36 ;
  END
END MUX2X4H7R

MACRO MUX2X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2X6H7R 0 0 ;
  SIZE 5.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.2 1.48 ;
        RECT 4.682 1.075 4.822 1.48 ;
        RECT 4.182 1.075 4.322 1.48 ;
        RECT 3.185 1.24 3.325 1.48 ;
        RECT 0.82 1.215 0.96 1.48 ;
        RECT 0.32 1.035 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.2 0.08 ;
        RECT 4.682 -0.08 4.822 0.326 ;
        RECT 4.182 -0.08 4.322 0.325 ;
        RECT 3.185 -0.08 3.325 0.16 ;
        RECT 0.82 -0.08 0.96 0.16 ;
        RECT 0.32 -0.08 0.41 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.72 0.655 1.06 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.06 0.655 3.4 0.745 ;
      LAYER MET2 ;
        RECT 3.25 0.43 3.35 0.96 ;
      LAYER VIA1 ;
        RECT 3.255 0.655 3.345 0.745 ;
    END
  END B
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.225 0.78 1.435 0.87 ;
        RECT 0.225 0.855 1.263 0.889 ;
        RECT 1.15 0.836 1.435 0.87 ;
        RECT 1.188 0.798 1.225 0.927 ;
        RECT 0.225 0.855 1.188 0.945 ;
        RECT 0.225 0.725 0.315 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.957 0.895 5.047 1.04 ;
        RECT 3.957 0.416 5.047 0.506 ;
        RECT 4.957 0.3 5.047 0.506 ;
        RECT 3.957 0.895 5.047 0.985 ;
        RECT 4.855 0.416 4.945 0.985 ;
        RECT 4.457 0.895 4.547 1.04 ;
        RECT 4.457 0.315 4.547 0.506 ;
        RECT 3.957 0.895 4.047 1.04 ;
        RECT 3.957 0.3 4.047 0.506 ;
      LAYER MET2 ;
        RECT 4.85 0.43 4.95 0.96 ;
      LAYER VIA1 ;
        RECT 4.855 0.655 4.945 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.38 1.14 3.066 1.23 ;
      RECT 1.38 1.14 3.108 1.209 ;
      RECT 1.38 1.14 3.146 1.169 ;
      RECT 3.777 0.17 3.867 1.15 ;
      RECT 3.028 1.121 3.867 1.15 ;
      RECT 3.108 1.06 3.867 1.15 ;
      RECT 3.066 1.081 3.867 1.15 ;
      RECT 3.777 0.655 4.574 0.745 ;
      RECT 3.107 0.25 3.401 0.34 ;
      RECT 3.065 0.25 3.443 0.319 ;
      RECT 3.027 0.25 3.481 0.279 ;
      RECT 3.443 0.17 3.867 0.26 ;
      RECT 3.363 0.231 3.867 0.26 ;
      RECT 3.401 0.191 3.443 0.319 ;
      RECT 1.38 0.231 3.145 0.26 ;
      RECT 1.38 0.191 3.107 0.26 ;
      RECT 1.38 0.17 3.065 0.26 ;
      RECT 2.345 0.92 3.015 1.01 ;
      RECT 2.925 0.88 3.605 0.97 ;
      RECT 3.515 0.43 3.605 0.97 ;
      RECT 2.912 0.43 3.687 0.52 ;
      RECT 3.547 0.355 3.687 0.52 ;
      RECT 2.87 0.371 2.912 0.499 ;
      RECT 2.832 0.43 3.687 0.459 ;
      RECT 1.935 0.35 2.87 0.44 ;
      RECT 1.935 0.411 2.95 0.44 ;
      RECT 0.54 1.035 1.265 1.125 ;
      RECT 0.54 1.035 1.302 1.107 ;
      RECT 0.54 1.035 1.34 1.069 ;
      RECT 2.165 0.53 2.255 1.05 ;
      RECT 1.227 1.016 2.255 1.05 ;
      RECT 1.302 0.96 2.255 1.05 ;
      RECT 1.265 0.978 2.255 1.05 ;
      RECT 1.725 0.53 2.255 0.62 ;
      RECT 1.725 0.35 1.815 0.62 ;
      RECT 1.302 0.35 1.815 0.44 ;
      RECT 1.286 0.304 1.302 0.432 ;
      RECT 1.24 0.273 1.286 0.401 ;
      RECT 1.202 0.331 1.34 0.359 ;
      RECT 0.54 0.25 1.24 0.34 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 0.045 0.28 0.135 1.13 ;
      RECT 1.661 0.74 2.075 0.83 ;
      RECT 1.627 0.685 1.661 0.813 ;
      RECT 1.581 0.645 1.627 0.773 ;
      RECT 1.581 0.721 1.699 0.773 ;
      RECT 1.535 0.599 1.581 0.727 ;
      RECT 1.489 0.553 1.535 0.681 ;
      RECT 1.451 0.599 1.581 0.639 ;
      RECT 1.225 0.53 1.489 0.62 ;
      RECT 1.208 0.483 1.225 0.612 ;
      RECT 1.17 0.553 1.535 0.584 ;
      RECT 0.045 0.475 1.208 0.565 ;
      RECT 0.045 0.511 1.263 0.565 ;
      RECT 0.045 0.28 0.185 0.37 ;
  END
END MUX2X6H7R

MACRO MUX2X8H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2X8H7R 0 0 ;
  SIZE 5.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.6 1.48 ;
        RECT 5.375 1.035 5.465 1.48 ;
        RECT 4.85 1.075 4.99 1.48 ;
        RECT 4.35 1.075 4.49 1.48 ;
        RECT 3.435 1.24 3.575 1.48 ;
        RECT 1.07 1.215 1.21 1.48 ;
        RECT 0.57 1.035 0.66 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.6 0.08 ;
        RECT 5.384 -0.08 5.474 0.359 ;
        RECT 4.859 -0.08 4.999 0.326 ;
        RECT 4.359 -0.08 4.499 0.325 ;
        RECT 3.362 -0.08 3.502 0.16 ;
        RECT 1.07 -0.08 1.21 0.205 ;
        RECT 0.585 -0.08 0.675 0.345 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.97 0.655 1.31 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.235 0.655 3.575 0.745 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END B
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.466 0.74 1.871 0.83 ;
        RECT 1.351 0.836 1.466 0.884 ;
        RECT 1.389 0.794 1.504 0.849 ;
        RECT 1.435 0.755 1.466 0.884 ;
        RECT 0.475 0.855 1.435 0.922 ;
        RECT 0.475 0.855 1.389 0.945 ;
        RECT 0.475 0.725 0.565 0.945 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.134 0.416 5.224 0.506 ;
        RECT 5.134 0.324 5.224 0.506 ;
        RECT 5.125 0.895 5.215 1.04 ;
        RECT 5.055 0.416 5.145 0.985 ;
        RECT 4.125 0.895 5.215 0.985 ;
        RECT 4.634 0.324 4.724 0.506 ;
        RECT 4.134 0.309 4.224 0.506 ;
        RECT 4.125 0.895 4.215 1.04 ;
      LAYER MET2 ;
        RECT 5.05 0.43 5.15 0.96 ;
      LAYER VIA1 ;
        RECT 5.055 0.655 5.145 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.705 1.139 3.317 1.229 ;
      RECT 1.705 1.139 3.358 1.209 ;
      RECT 1.705 1.139 3.396 1.169 ;
      RECT 3.945 0.17 4.035 1.15 ;
      RECT 3.279 1.12 4.035 1.15 ;
      RECT 3.358 1.06 4.035 1.15 ;
      RECT 3.317 1.08 4.035 1.15 ;
      RECT 3.945 0.655 4.824 0.745 ;
      RECT 3.284 0.25 3.584 0.34 ;
      RECT 3.242 0.25 3.626 0.319 ;
      RECT 3.204 0.25 3.664 0.279 ;
      RECT 3.626 0.17 4.035 0.26 ;
      RECT 3.546 0.231 4.035 0.26 ;
      RECT 3.584 0.191 3.626 0.319 ;
      RECT 1.63 0.231 3.322 0.26 ;
      RECT 1.63 0.191 3.284 0.26 ;
      RECT 1.63 0.17 3.242 0.26 ;
      RECT 2.595 0.9 3.265 0.99 ;
      RECT 3.765 0.35 3.855 0.97 ;
      RECT 3.175 0.88 3.855 0.97 ;
      RECT 3.162 0.43 3.855 0.52 ;
      RECT 3.715 0.35 3.855 0.52 ;
      RECT 3.12 0.371 3.162 0.499 ;
      RECT 3.082 0.43 3.855 0.459 ;
      RECT 2.213 0.35 3.12 0.44 ;
      RECT 2.213 0.411 3.2 0.44 ;
      RECT 0.79 1.035 1.515 1.125 ;
      RECT 0.79 1.035 1.553 1.106 ;
      RECT 0.79 1.035 1.591 1.068 ;
      RECT 2.415 0.53 2.505 1.049 ;
      RECT 1.477 1.016 2.505 1.049 ;
      RECT 1.553 0.959 2.505 1.049 ;
      RECT 1.515 0.978 2.505 1.049 ;
      RECT 2.137 0.53 2.505 0.62 ;
      RECT 2.127 0.487 2.137 0.615 ;
      RECT 2.081 0.459 2.127 0.587 ;
      RECT 2.035 0.413 2.081 0.541 ;
      RECT 2.035 0.511 2.175 0.541 ;
      RECT 2.003 0.35 2.035 0.502 ;
      RECT 1.957 0.35 2.035 0.463 ;
      RECT 1.552 0.35 2.035 0.44 ;
      RECT 1.535 0.303 1.552 0.432 ;
      RECT 1.497 0.35 2.035 0.404 ;
      RECT 0.79 0.295 1.535 0.385 ;
      RECT 0.79 0.331 1.59 0.385 ;
      RECT 0.295 1.03 0.435 1.12 ;
      RECT 0.295 0.245 0.385 1.12 ;
      RECT 2.215 0.715 2.305 0.855 ;
      RECT 2.066 0.715 2.305 0.805 ;
      RECT 2.062 0.675 2.066 0.803 ;
      RECT 2.016 0.65 2.062 0.778 ;
      RECT 1.97 0.604 2.016 0.732 ;
      RECT 1.97 0.696 2.104 0.732 ;
      RECT 1.924 0.558 1.97 0.686 ;
      RECT 1.886 0.604 2.016 0.644 ;
      RECT 1.45 0.535 1.924 0.625 ;
      RECT 1.428 0.486 1.45 0.614 ;
      RECT 1.39 0.558 1.97 0.584 ;
      RECT 0.295 0.475 1.428 0.565 ;
      RECT 0.295 0.516 1.488 0.565 ;
      RECT 0.295 0.245 0.435 0.335 ;
  END
END MUX2X8H7R

MACRO MUX4X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX4X0P5H7R 0 0 ;
  SIZE 4.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.6 1.48 ;
        RECT 4.035 0.959 4.125 1.48 ;
        RECT 2.322 1.095 2.462 1.48 ;
        RECT 1.53 1.07 1.62 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.6 0.08 ;
        RECT 4.045 -0.08 4.135 0.33 ;
        RECT 2.527 -0.08 2.617 0.38 ;
        RECT 1.515 -0.08 1.605 0.38 ;
        RECT 0.295 -0.08 0.435 0.342 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.355 0.655 2.58 0.775 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.605 0.65 1.875 0.75 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.655 0.59 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.215 0.655 1.515 0.745 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END D
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.71 0.455 0.8 0.845 ;
        RECT 0.225 0.455 0.8 0.545 ;
        RECT 0.225 0.455 0.315 0.61 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END S0
  PIN S1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.875 0.455 4.175 0.545 ;
      LAYER MET2 ;
        RECT 4.05 0.23 4.15 0.76 ;
      LAYER VIA1 ;
        RECT 4.055 0.455 4.145 0.545 ;
    END
  END S1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.315 0.205 4.405 1.044 ;
        RECT 4.225 0.205 4.405 0.345 ;
      LAYER MET2 ;
        RECT 4.25 0.18 4.35 0.56 ;
      LAYER VIA1 ;
        RECT 4.255 0.255 4.345 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 3.182 1.14 3.937 1.23 ;
      RECT 3.847 0.862 3.937 1.23 ;
      RECT 3.182 0.35 3.272 1.23 ;
      RECT 3.847 0.862 3.983 0.9 ;
      RECT 3.893 0.817 3.988 0.875 ;
      RECT 3.893 0.817 4.026 0.853 ;
      RECT 4.135 0.694 4.225 0.834 ;
      RECT 3.937 0.772 4.225 0.834 ;
      RECT 3.988 0.744 4.225 0.834 ;
      RECT 3.983 0.746 4.225 0.834 ;
      RECT 3.182 0.35 3.337 0.44 ;
      RECT 3.667 0.645 3.757 1.045 ;
      RECT 3.682 0.23 3.772 0.735 ;
      RECT 3.682 0.23 3.91 0.32 ;
      RECT 0.869 0.96 1.009 1.05 ;
      RECT 0.919 0.445 1.009 1.05 ;
      RECT 3.407 0.86 3.577 0.95 ;
      RECT 3.487 0.469 3.577 0.95 ;
      RECT 2.347 0.47 2.797 0.56 ;
      RECT 2.707 0.17 2.797 0.56 ;
      RECT 1.335 0.47 1.785 0.56 ;
      RECT 1.695 0.265 1.785 0.56 ;
      RECT 0.919 0.445 1.425 0.535 ;
      RECT 3.502 0.17 3.592 0.508 ;
      RECT 2.347 0.265 2.437 0.56 ;
      RECT 1.695 0.265 2.437 0.355 ;
      RECT 2.707 0.17 3.592 0.26 ;
      RECT 2.102 0.445 2.192 1.155 ;
      RECT 2.807 0.915 2.897 1.14 ;
      RECT 2.102 0.915 2.977 1.005 ;
      RECT 2.887 0.35 2.977 1.005 ;
      RECT 1.965 0.445 2.192 0.535 ;
      RECT 2.887 0.35 3.027 0.44 ;
      RECT 0.578 1.14 1.205 1.23 ;
      RECT 1.115 0.841 1.205 1.23 ;
      RECT 0.045 0.915 0.16 1.155 ;
      RECT 0.578 1.028 0.668 1.23 ;
      RECT 0.533 0.937 0.578 1.066 ;
      RECT 0.533 0.983 0.624 1.066 ;
      RECT 0.495 0.983 0.624 1.024 ;
      RECT 0.045 0.915 0.533 1.005 ;
      RECT 1.115 0.841 2.012 0.931 ;
      RECT 0.045 0.267 0.135 1.155 ;
      RECT 0.045 0.267 0.185 0.357 ;
  END
END MUX4X0P5H7R

MACRO MUX4X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX4X0P7H7R 0 0 ;
  SIZE 4.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.6 1.48 ;
        RECT 4.035 0.991 4.125 1.48 ;
        RECT 2.322 1.095 2.462 1.48 ;
        RECT 1.53 1.07 1.62 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.6 0.08 ;
        RECT 4.045 -0.08 4.135 0.33 ;
        RECT 2.527 -0.08 2.617 0.38 ;
        RECT 1.515 -0.08 1.605 0.38 ;
        RECT 0.295 -0.08 0.435 0.342 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.355 0.655 2.58 0.775 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.605 0.65 1.875 0.75 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.655 0.59 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.215 0.655 1.515 0.745 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END D
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.71 0.455 0.8 0.845 ;
        RECT 0.225 0.455 0.8 0.545 ;
        RECT 0.225 0.455 0.315 0.61 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END S0
  PIN S1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.875 0.455 4.175 0.545 ;
      LAYER MET2 ;
        RECT 4.05 0.23 4.15 0.76 ;
      LAYER VIA1 ;
        RECT 4.055 0.455 4.145 0.545 ;
    END
  END S1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.315 0.229 4.405 1.044 ;
        RECT 4.225 0.229 4.405 0.36 ;
      LAYER MET2 ;
        RECT 4.25 0.18 4.35 0.56 ;
      LAYER VIA1 ;
        RECT 4.255 0.255 4.345 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 3.182 1.14 3.937 1.23 ;
      RECT 3.847 0.862 3.937 1.23 ;
      RECT 3.182 0.35 3.272 1.23 ;
      RECT 3.847 0.862 3.983 0.9 ;
      RECT 3.893 0.817 3.988 0.875 ;
      RECT 3.893 0.817 4.026 0.853 ;
      RECT 4.135 0.694 4.225 0.834 ;
      RECT 3.937 0.772 4.225 0.834 ;
      RECT 3.988 0.744 4.225 0.834 ;
      RECT 3.983 0.746 4.225 0.834 ;
      RECT 3.182 0.35 3.337 0.44 ;
      RECT 3.667 0.645 3.757 1.045 ;
      RECT 3.682 0.23 3.772 0.695 ;
      RECT 3.682 0.23 3.91 0.32 ;
      RECT 0.869 0.96 1.009 1.05 ;
      RECT 0.919 0.445 1.009 1.05 ;
      RECT 3.407 0.86 3.577 0.95 ;
      RECT 3.487 0.469 3.577 0.95 ;
      RECT 2.347 0.47 2.797 0.56 ;
      RECT 2.707 0.17 2.797 0.56 ;
      RECT 1.335 0.47 1.785 0.56 ;
      RECT 1.695 0.265 1.785 0.56 ;
      RECT 0.919 0.445 1.425 0.535 ;
      RECT 3.502 0.17 3.592 0.508 ;
      RECT 2.347 0.265 2.437 0.56 ;
      RECT 1.695 0.265 2.437 0.355 ;
      RECT 2.707 0.17 3.592 0.26 ;
      RECT 2.102 0.445 2.192 1.155 ;
      RECT 2.807 0.915 2.897 1.14 ;
      RECT 2.102 0.915 2.977 1.005 ;
      RECT 2.887 0.35 2.977 1.005 ;
      RECT 1.965 0.445 2.192 0.535 ;
      RECT 2.887 0.35 3.027 0.44 ;
      RECT 0.578 1.14 1.205 1.23 ;
      RECT 1.115 0.841 1.205 1.23 ;
      RECT 0.045 0.915 0.16 1.155 ;
      RECT 0.578 1.028 0.668 1.23 ;
      RECT 0.533 0.937 0.578 1.066 ;
      RECT 0.533 0.983 0.624 1.066 ;
      RECT 0.495 0.983 0.624 1.024 ;
      RECT 0.045 0.915 0.533 1.005 ;
      RECT 1.115 0.841 2.012 0.931 ;
      RECT 0.045 0.267 0.135 1.155 ;
      RECT 0.045 0.267 0.185 0.357 ;
  END
END MUX4X0P7H7R

MACRO MUX4X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX4X1H7R 0 0 ;
  SIZE 4.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.6 1.48 ;
        RECT 4.035 1.039 4.125 1.48 ;
        RECT 2.322 1.095 2.462 1.48 ;
        RECT 1.53 1.07 1.62 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.6 0.08 ;
        RECT 4.045 -0.08 4.135 0.33 ;
        RECT 2.527 -0.08 2.617 0.38 ;
        RECT 1.515 -0.08 1.605 0.38 ;
        RECT 0.295 -0.08 0.435 0.342 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.355 0.655 2.58 0.775 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.605 0.65 1.875 0.75 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.655 0.59 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.215 0.655 1.515 0.745 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END D
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.71 0.455 0.8 0.845 ;
        RECT 0.225 0.455 0.8 0.545 ;
        RECT 0.225 0.455 0.315 0.61 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END S0
  PIN S1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.875 0.455 4.175 0.545 ;
      LAYER MET2 ;
        RECT 4.05 0.23 4.15 0.76 ;
      LAYER VIA1 ;
        RECT 4.055 0.455 4.145 0.545 ;
    END
  END S1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.315 0.255 4.405 1.044 ;
        RECT 4.225 0.255 4.405 0.345 ;
      LAYER MET2 ;
        RECT 4.25 0.18 4.35 0.56 ;
      LAYER VIA1 ;
        RECT 4.255 0.255 4.345 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 3.182 1.14 3.937 1.23 ;
      RECT 3.847 0.862 3.937 1.23 ;
      RECT 3.182 0.35 3.272 1.23 ;
      RECT 3.847 0.862 3.983 0.9 ;
      RECT 3.893 0.817 3.988 0.875 ;
      RECT 3.893 0.817 4.026 0.853 ;
      RECT 4.135 0.694 4.225 0.834 ;
      RECT 3.937 0.772 4.225 0.834 ;
      RECT 3.988 0.744 4.225 0.834 ;
      RECT 3.983 0.746 4.225 0.834 ;
      RECT 3.182 0.35 3.337 0.44 ;
      RECT 3.667 0.645 3.757 1.045 ;
      RECT 3.682 0.23 3.772 0.735 ;
      RECT 3.682 0.23 3.91 0.32 ;
      RECT 0.869 0.96 1.009 1.05 ;
      RECT 0.919 0.445 1.009 1.05 ;
      RECT 3.407 0.86 3.577 0.95 ;
      RECT 3.487 0.469 3.577 0.95 ;
      RECT 2.347 0.47 2.797 0.56 ;
      RECT 2.707 0.17 2.797 0.56 ;
      RECT 1.335 0.47 1.785 0.56 ;
      RECT 1.695 0.265 1.785 0.56 ;
      RECT 0.919 0.445 1.425 0.535 ;
      RECT 3.502 0.17 3.592 0.508 ;
      RECT 2.347 0.265 2.437 0.56 ;
      RECT 1.695 0.265 2.437 0.355 ;
      RECT 2.707 0.17 3.592 0.26 ;
      RECT 2.102 0.445 2.192 1.155 ;
      RECT 2.807 0.915 2.897 1.14 ;
      RECT 2.102 0.915 2.977 1.005 ;
      RECT 2.887 0.35 2.977 1.005 ;
      RECT 1.965 0.445 2.192 0.535 ;
      RECT 2.887 0.35 3.027 0.44 ;
      RECT 0.578 1.14 1.205 1.23 ;
      RECT 1.115 0.841 1.205 1.23 ;
      RECT 0.045 0.915 0.16 1.155 ;
      RECT 0.578 1.028 0.668 1.23 ;
      RECT 0.533 0.937 0.578 1.066 ;
      RECT 0.533 0.983 0.624 1.066 ;
      RECT 0.495 0.983 0.624 1.024 ;
      RECT 0.045 0.915 0.533 1.005 ;
      RECT 1.115 0.841 2.012 0.931 ;
      RECT 0.045 0.267 0.135 1.155 ;
      RECT 0.045 0.267 0.185 0.357 ;
  END
END MUX4X1H7R

MACRO MUX4X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX4X1P4H7R 0 0 ;
  SIZE 4.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.6 1.48 ;
        RECT 4.035 1.07 4.125 1.48 ;
        RECT 2.322 1.095 2.462 1.48 ;
        RECT 1.53 1.07 1.62 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.6 0.08 ;
        RECT 4.045 -0.08 4.135 0.33 ;
        RECT 2.527 -0.08 2.617 0.38 ;
        RECT 1.515 -0.08 1.605 0.38 ;
        RECT 0.295 -0.08 0.435 0.342 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.39 0.65 2.59 0.785 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.605 0.65 1.875 0.75 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.655 0.59 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.215 0.655 1.515 0.745 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END D
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.71 0.455 0.8 0.845 ;
        RECT 0.225 0.455 0.8 0.545 ;
        RECT 0.225 0.455 0.315 0.61 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END S0
  PIN S1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.885 0.455 4.175 0.55 ;
      LAYER MET2 ;
        RECT 4.05 0.23 4.15 0.76 ;
      LAYER VIA1 ;
        RECT 4.055 0.455 4.145 0.545 ;
    END
  END S1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.315 0.255 4.405 1.031 ;
        RECT 4.225 0.255 4.405 0.345 ;
      LAYER MET2 ;
        RECT 4.25 0.18 4.35 0.56 ;
      LAYER VIA1 ;
        RECT 4.255 0.255 4.345 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 3.182 1.14 3.937 1.23 ;
      RECT 3.847 0.755 3.937 1.23 ;
      RECT 3.182 0.35 3.272 1.23 ;
      RECT 3.847 0.755 4.225 0.845 ;
      RECT 4.135 0.705 4.225 0.845 ;
      RECT 3.182 0.35 3.337 0.44 ;
      RECT 3.667 0.371 3.757 1.035 ;
      RECT 3.713 0.326 3.816 0.396 ;
      RECT 3.757 0.297 3.77 0.426 ;
      RECT 3.77 0.23 3.862 0.35 ;
      RECT 3.757 0.297 3.869 0.324 ;
      RECT 3.77 0.23 3.91 0.32 ;
      RECT 0.869 0.96 1.009 1.05 ;
      RECT 0.919 0.445 1.009 1.05 ;
      RECT 3.407 0.86 3.577 0.95 ;
      RECT 3.487 0.17 3.577 0.95 ;
      RECT 2.347 0.47 2.797 0.56 ;
      RECT 2.707 0.17 2.797 0.56 ;
      RECT 1.335 0.47 1.785 0.56 ;
      RECT 1.695 0.17 1.785 0.56 ;
      RECT 0.919 0.445 1.425 0.535 ;
      RECT 2.347 0.17 2.437 0.56 ;
      RECT 3.487 0.17 3.592 0.33 ;
      RECT 2.707 0.17 3.592 0.26 ;
      RECT 1.695 0.17 2.437 0.26 ;
      RECT 2.102 0.445 2.192 1.155 ;
      RECT 2.807 0.915 2.897 1.14 ;
      RECT 2.102 0.915 2.977 1.005 ;
      RECT 2.887 0.36 2.977 1.005 ;
      RECT 1.965 0.445 2.192 0.535 ;
      RECT 2.887 0.36 3.027 0.45 ;
      RECT 0.578 1.14 1.205 1.23 ;
      RECT 1.115 0.841 1.205 1.23 ;
      RECT 0.045 0.915 0.16 1.155 ;
      RECT 0.578 1.028 0.668 1.23 ;
      RECT 0.533 0.937 0.578 1.066 ;
      RECT 0.533 0.983 0.624 1.066 ;
      RECT 0.495 0.983 0.624 1.024 ;
      RECT 0.045 0.915 0.533 1.005 ;
      RECT 1.115 0.841 2.012 0.931 ;
      RECT 0.045 0.242 0.135 1.155 ;
      RECT 0.045 0.242 0.16 0.382 ;
  END
END MUX4X1P4H7R

MACRO MUX4X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX4X2H7R 0 0 ;
  SIZE 4.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.8 1.48 ;
        RECT 4.53 0.945 4.62 1.48 ;
        RECT 4.03 0.959 4.12 1.48 ;
        RECT 2.322 1.095 2.462 1.48 ;
        RECT 1.53 1.07 1.62 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.8 0.08 ;
        RECT 4.53 -0.08 4.62 0.345 ;
        RECT 3.992 -0.08 4.082 0.33 ;
        RECT 2.527 -0.08 2.617 0.38 ;
        RECT 1.515 -0.08 1.605 0.38 ;
        RECT 0.295 -0.08 0.435 0.342 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.402 0.65 2.602 0.785 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.605 0.65 1.875 0.75 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.655 0.59 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.215 0.655 1.515 0.745 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END D
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.71 0.455 0.8 0.845 ;
        RECT 0.225 0.455 0.8 0.545 ;
        RECT 0.225 0.455 0.315 0.61 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END S0
  PIN S1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.857 0.455 4.175 0.545 ;
      LAYER MET2 ;
        RECT 4.05 0.23 4.15 0.76 ;
      LAYER VIA1 ;
        RECT 4.055 0.455 4.145 0.545 ;
    END
  END S1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.255 0.915 4.4 1.005 ;
        RECT 4.31 0.245 4.4 1.005 ;
        RECT 4.217 0.245 4.4 0.345 ;
      LAYER MET2 ;
        RECT 4.25 0.18 4.35 0.56 ;
      LAYER VIA1 ;
        RECT 4.255 0.255 4.345 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 3.182 1.14 3.932 1.23 ;
      RECT 3.842 0.735 3.932 1.23 ;
      RECT 3.182 0.35 3.272 1.23 ;
      RECT 3.842 0.735 4.22 0.825 ;
      RECT 4.13 0.685 4.22 0.825 ;
      RECT 3.182 0.35 3.337 0.44 ;
      RECT 3.662 0.371 3.752 1.05 ;
      RECT 3.708 0.331 3.798 0.409 ;
      RECT 3.742 0.205 3.832 0.369 ;
      RECT 0.869 0.96 1.009 1.05 ;
      RECT 0.919 0.445 1.009 1.05 ;
      RECT 3.407 0.86 3.572 0.95 ;
      RECT 3.482 0.17 3.572 0.95 ;
      RECT 2.347 0.47 2.797 0.56 ;
      RECT 2.707 0.17 2.797 0.56 ;
      RECT 1.335 0.47 1.785 0.56 ;
      RECT 1.695 0.265 1.785 0.56 ;
      RECT 0.919 0.445 1.425 0.535 ;
      RECT 2.347 0.265 2.437 0.56 ;
      RECT 1.695 0.265 2.437 0.355 ;
      RECT 3.482 0.17 3.592 0.34 ;
      RECT 2.707 0.17 3.592 0.26 ;
      RECT 2.102 0.445 2.192 1.163 ;
      RECT 2.807 0.915 2.897 1.14 ;
      RECT 2.102 0.915 2.977 1.005 ;
      RECT 2.887 0.35 2.977 1.005 ;
      RECT 1.965 0.445 2.192 0.535 ;
      RECT 2.887 0.35 3.027 0.44 ;
      RECT 0.578 1.14 1.205 1.23 ;
      RECT 1.115 0.841 1.205 1.23 ;
      RECT 0.045 0.915 0.16 1.155 ;
      RECT 0.578 1.028 0.668 1.23 ;
      RECT 0.533 0.937 0.578 1.066 ;
      RECT 0.533 0.983 0.624 1.066 ;
      RECT 0.495 0.983 0.624 1.024 ;
      RECT 0.045 0.915 0.533 1.005 ;
      RECT 1.115 0.841 2.012 0.931 ;
      RECT 0.045 0.242 0.135 1.155 ;
      RECT 0.045 0.242 0.16 0.382 ;
  END
END MUX4X2H7R

MACRO MUX4X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX4X3H7R 0 0 ;
  SIZE 5 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5 1.48 ;
        RECT 4.719 1.04 4.809 1.48 ;
        RECT 4.219 1.055 4.309 1.48 ;
        RECT 2.531 1.055 2.621 1.48 ;
        RECT 1.608 1.07 1.698 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5 0.08 ;
        RECT 4.719 -0.08 4.809 0.345 ;
        RECT 4.181 -0.08 4.271 0.33 ;
        RECT 2.711 -0.08 2.801 0.38 ;
        RECT 1.571 -0.08 1.711 0.325 ;
        RECT 0.295 -0.08 0.435 0.342 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.586 0.65 2.786 0.785 ;
      LAYER MET2 ;
        RECT 2.65 0.43 2.75 0.96 ;
      LAYER VIA1 ;
        RECT 2.655 0.655 2.745 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.715 0.655 1.975 0.78 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.405 0.655 0.585 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.396 0.645 1.596 0.78 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END D
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.705 0.455 0.795 0.845 ;
        RECT 0.225 0.455 0.795 0.545 ;
        RECT 0.225 0.455 0.315 0.642 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END S0
  PIN S1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.051 0.495 4.345 0.585 ;
        RECT 4.255 0.425 4.345 0.585 ;
      LAYER MET2 ;
        RECT 4.25 0.225 4.35 0.76 ;
      LAYER VIA1 ;
        RECT 4.255 0.455 4.345 0.545 ;
    END
  END S1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.444 0.94 4.623 1.03 ;
        RECT 4.533 0.255 4.623 1.03 ;
        RECT 4.406 0.255 4.623 0.345 ;
      LAYER MET2 ;
        RECT 4.45 0.18 4.55 0.56 ;
      LAYER VIA1 ;
        RECT 4.455 0.255 4.545 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 3.351 1.14 4.121 1.23 ;
      RECT 4.031 0.849 4.121 1.23 ;
      RECT 3.351 0.35 3.441 1.23 ;
      RECT 4.077 0.804 4.186 0.864 ;
      RECT 4.121 0.768 4.148 0.897 ;
      RECT 4.319 0.705 4.409 0.845 ;
      RECT 4.148 0.755 4.409 0.845 ;
      RECT 3.351 0.35 3.491 0.44 ;
      RECT 3.851 0.38 3.941 1.05 ;
      RECT 3.897 0.34 3.987 0.418 ;
      RECT 3.931 0.205 4.021 0.378 ;
      RECT 0.795 0.96 1.031 1.05 ;
      RECT 0.941 0.415 1.031 1.05 ;
      RECT 3.591 0.86 3.761 0.95 ;
      RECT 3.671 0.17 3.761 0.95 ;
      RECT 2.531 0.47 2.981 0.56 ;
      RECT 2.891 0.17 2.981 0.56 ;
      RECT 0.941 0.415 1.891 0.505 ;
      RECT 1.801 0.265 1.891 0.505 ;
      RECT 2.531 0.265 2.621 0.56 ;
      RECT 1.801 0.265 2.621 0.355 ;
      RECT 3.671 0.17 3.781 0.345 ;
      RECT 2.891 0.17 3.781 0.26 ;
      RECT 2.155 1.05 2.441 1.14 ;
      RECT 2.351 0.445 2.441 1.14 ;
      RECT 2.991 0.875 3.081 1.08 ;
      RECT 2.351 0.875 3.161 0.965 ;
      RECT 3.071 0.35 3.161 0.965 ;
      RECT 2.046 0.445 2.441 0.535 ;
      RECT 3.071 0.35 3.211 0.44 ;
      RECT 0.578 1.14 1.311 1.23 ;
      RECT 1.221 0.87 1.311 1.23 ;
      RECT 0.045 0.915 0.16 1.155 ;
      RECT 0.578 1.04 0.668 1.23 ;
      RECT 0.567 0.966 0.578 1.095 ;
      RECT 0.521 0.938 0.567 1.066 ;
      RECT 0.521 0.995 0.624 1.066 ;
      RECT 0.483 0.995 0.624 1.024 ;
      RECT 0.045 0.915 0.521 1.005 ;
      RECT 1.221 0.87 2.261 0.96 ;
      RECT 2.171 0.736 2.261 0.96 ;
      RECT 0.045 0.242 0.135 1.155 ;
      RECT 0.045 0.242 0.16 0.382 ;
  END
END MUX4X3H7R

MACRO MUX4X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX4X4H7R 0 0 ;
  SIZE 5.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.8 1.48 ;
        RECT 5.39 1.045 5.48 1.48 ;
        RECT 4.89 1.045 4.98 1.48 ;
        RECT 3.268 1.03 3.358 1.48 ;
        RECT 1.958 1.24 2.098 1.48 ;
        RECT 0.795 1.24 0.935 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.8 0.08 ;
        RECT 5.378 -0.08 5.468 0.33 ;
        RECT 4.855 -0.08 4.945 0.33 ;
        RECT 3.354 -0.08 3.494 0.16 ;
        RECT 1.908 -0.08 2.048 0.16 ;
        RECT 0.795 -0.08 0.935 0.16 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.245 0.625 3.425 0.775 ;
      LAYER MET2 ;
        RECT 3.25 0.43 3.35 0.96 ;
      LAYER VIA1 ;
        RECT 3.255 0.655 3.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.025 0.455 2.2 0.61 ;
      LAYER MET2 ;
        RECT 2.05 0.23 2.15 0.76 ;
      LAYER VIA1 ;
        RECT 2.055 0.455 2.145 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.64 0.625 0.82 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.975 0.625 1.155 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END D
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.588 0.89 2.973 0.98 ;
        RECT 2.883 0.66 2.973 0.98 ;
        RECT 1.803 0.7 2.973 0.79 ;
        RECT 1.598 1.06 2.678 1.15 ;
        RECT 2.588 0.89 2.678 1.15 ;
        RECT 2.373 0.51 2.463 0.79 ;
        RECT 1.803 0.645 1.893 0.79 ;
        RECT 1.502 1.041 1.636 1.077 ;
        RECT 1.502 1.02 1.598 1.077 ;
        RECT 1.594 1.06 2.678 1.148 ;
        RECT 1.456 0.995 1.594 1.031 ;
        RECT 1.548 1.06 2.678 1.123 ;
        RECT 1.456 0.949 1.548 1.031 ;
        RECT 0.425 0.903 1.502 0.97 ;
        RECT 0.425 0.88 1.456 0.97 ;
        RECT 1.418 0.949 1.548 0.989 ;
        RECT 0.425 0.855 0.575 0.97 ;
        RECT 0.455 0.665 0.545 0.97 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END S0
  PIN S1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.765 0.455 4.975 0.595 ;
      LAYER MET2 ;
        RECT 4.85 0.23 4.95 0.76 ;
      LAYER VIA1 ;
        RECT 4.855 0.455 4.945 0.545 ;
    END
  END S1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.64 0.255 5.73 1.08 ;
        RECT 5.198 0.655 5.73 0.745 ;
        RECT 5.115 0.955 5.288 1.045 ;
        RECT 5.198 0.295 5.288 1.045 ;
        RECT 5.08 0.295 5.288 0.385 ;
      LAYER MET2 ;
        RECT 5.45 0.425 5.55 0.96 ;
      LAYER VIA1 ;
        RECT 5.455 0.655 5.545 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 3.795 1.11 4.8 1.2 ;
      RECT 4.71 0.72 4.8 1.2 ;
      RECT 4.295 0.855 4.385 1.2 ;
      RECT 3.795 0.637 3.885 1.2 ;
      RECT 4.71 0.72 5.108 0.81 ;
      RECT 3.795 0.637 3.931 0.675 ;
      RECT 3.841 0.592 3.94 0.648 ;
      RECT 3.885 0.547 3.986 0.62 ;
      RECT 3.931 0.519 3.94 0.648 ;
      RECT 3.94 0.35 4.03 0.575 ;
      RECT 3.94 0.35 4.08 0.44 ;
      RECT 4.525 0.797 4.615 1.02 ;
      RECT 4.499 0.797 4.615 0.835 ;
      RECT 4.453 0.452 4.543 0.799 ;
      RECT 4.453 0.761 4.589 0.799 ;
      RECT 4.453 0.452 4.589 0.49 ;
      RECT 4.499 0.416 4.605 0.459 ;
      RECT 4.525 0.394 4.651 0.428 ;
      RECT 4.589 0.331 4.605 0.459 ;
      RECT 4.543 0.362 4.651 0.428 ;
      RECT 4.605 0.205 4.695 0.383 ;
      RECT 1.201 1.14 1.46 1.23 ;
      RECT 0.302 1.06 1.083 1.15 ;
      RECT 4.02 0.86 4.073 0.95 ;
      RECT 0.135 0.265 1.445 0.355 ;
      RECT 1.355 0.17 1.445 0.355 ;
      RECT 3.274 0.25 3.532 0.34 ;
      RECT 1.869 0.25 2.087 0.34 ;
      RECT 3.65 0.17 4.215 0.26 ;
      RECT 2.205 0.17 3.156 0.26 ;
      RECT 1.355 0.17 1.751 0.26 ;
      RECT 4.261 0.17 4.305 0.676 ;
      RECT 4.215 0.17 4.261 0.721 ;
      RECT 4.209 0.619 4.215 0.747 ;
      RECT 4.163 0.645 4.209 0.773 ;
      RECT 4.119 0.69 4.163 0.95 ;
      RECT 4.073 0.735 4.119 0.95 ;
      RECT 3.612 0.17 3.65 0.279 ;
      RECT 3.57 0.191 3.612 0.319 ;
      RECT 3.532 0.231 3.57 0.34 ;
      RECT 3.236 0.231 3.274 0.34 ;
      RECT 3.194 0.191 3.236 0.319 ;
      RECT 3.156 0.17 3.194 0.279 ;
      RECT 2.167 0.17 2.205 0.279 ;
      RECT 2.125 0.191 2.167 0.319 ;
      RECT 2.087 0.231 2.125 0.34 ;
      RECT 1.831 0.231 1.869 0.34 ;
      RECT 1.789 0.191 1.831 0.319 ;
      RECT 1.751 0.17 1.789 0.279 ;
      RECT 1.163 1.121 1.201 1.23 ;
      RECT 1.121 1.081 1.163 1.209 ;
      RECT 1.083 1.06 1.121 1.169 ;
      RECT 0.264 1.041 0.302 1.15 ;
      RECT 0.227 1.003 0.264 1.132 ;
      RECT 0.181 0.962 0.227 1.09 ;
      RECT 0.135 0.916 0.181 1.044 ;
      RECT 0.091 0.265 0.135 0.999 ;
      RECT 0.045 0.265 0.091 0.954 ;
      RECT 2.768 1.07 3.153 1.16 ;
      RECT 3.063 0.43 3.153 1.16 ;
      RECT 3.499 0.92 3.705 1.01 ;
      RECT 3.615 0.401 3.705 1.01 ;
      RECT 3.661 0.364 3.705 1.01 ;
      RECT 3.063 0.43 3.705 0.52 ;
      RECT 3.609 0.427 3.705 0.52 ;
      RECT 3.049 0.357 3.063 0.485 ;
      RECT 3.011 0.43 3.705 0.459 ;
      RECT 3.011 0.43 3.727 0.451 ;
      RECT 3.689 0.35 3.83 0.44 ;
      RECT 2.528 0.42 3.129 0.44 ;
      RECT 2.528 0.387 3.109 0.44 ;
      RECT 2.528 0.35 3.049 0.44 ;
      RECT 1.674 0.88 2.498 0.97 ;
      RECT 1.663 0.836 1.674 0.965 ;
      RECT 1.619 0.88 2.498 0.937 ;
      RECT 1.573 0.35 1.663 0.892 ;
      RECT 1.573 0.861 1.712 0.892 ;
      RECT 1.53 0.69 1.663 0.848 ;
      RECT 1.484 0.69 1.663 0.803 ;
      RECT 1.415 0.69 1.663 0.78 ;
      RECT 0.225 0.445 0.315 0.655 ;
      RECT 0.225 0.445 1.663 0.535 ;
      RECT 1.573 0.35 1.713 0.44 ;
  END
END MUX4X4H7R

MACRO MUX4X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX4X6H7R 0 0 ;
  SIZE 7 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7 1.48 ;
        RECT 6.766 1.055 6.856 1.48 ;
        RECT 6.241 1.095 6.381 1.48 ;
        RECT 5.766 1.015 5.856 1.48 ;
        RECT 4.141 1.055 4.231 1.48 ;
        RECT 2.636 1.24 2.776 1.48 ;
        RECT 1.112 1.24 1.252 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7 0.08 ;
        RECT 6.766 -0.08 6.856 0.345 ;
        RECT 6.266 -0.08 6.356 0.33 ;
        RECT 5.728 -0.08 5.818 0.33 ;
        RECT 4.196 -0.08 4.336 0.16 ;
        RECT 2.636 -0.08 2.776 0.16 ;
        RECT 1.112 -0.08 1.252 0.16 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.165 0.625 4.345 0.775 ;
      LAYER MET2 ;
        RECT 4.25 0.425 4.35 0.96 ;
      LAYER VIA1 ;
        RECT 4.255 0.655 4.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.625 0.445 2.79 0.61 ;
      LAYER MET2 ;
        RECT 2.65 0.23 2.75 0.76 ;
      LAYER VIA1 ;
        RECT 2.655 0.455 2.745 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.92 0.64 1.18 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.317 0.64 1.575 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END D
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.466 0.915 3.871 1.005 ;
        RECT 3.781 0.64 3.871 1.005 ;
        RECT 2.426 0.7 3.871 0.79 ;
        RECT 2.225 1.06 3.556 1.15 ;
        RECT 3.466 0.915 3.556 1.15 ;
        RECT 3.121 0.593 3.211 0.79 ;
        RECT 2.426 0.615 2.516 0.79 ;
        RECT 2.15 1.041 2.263 1.098 ;
        RECT 2.104 1.007 2.225 1.052 ;
        RECT 2.196 1.06 3.556 1.136 ;
        RECT 2.104 0.97 2.196 1.052 ;
        RECT 2.058 0.924 2.15 1.006 ;
        RECT 0.727 0.878 2.104 0.945 ;
        RECT 0.727 0.855 2.058 0.945 ;
        RECT 2.02 0.924 2.15 0.964 ;
        RECT 0.727 0.61 0.817 0.945 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END S0
  PIN S1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.6 0.455 5.78 0.605 ;
      LAYER MET2 ;
        RECT 5.65 0.225 5.75 0.76 ;
      LAYER VIA1 ;
        RECT 5.655 0.455 5.745 0.545 ;
    END
  END S1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.516 0.295 6.606 1.055 ;
        RECT 6.016 0.915 6.606 1.005 ;
        RECT 5.978 0.455 6.606 0.545 ;
        RECT 6.016 0.915 6.106 1.055 ;
        RECT 5.978 0.295 6.068 0.545 ;
      LAYER MET2 ;
        RECT 6.45 0.225 6.55 0.76 ;
      LAYER VIA1 ;
        RECT 6.455 0.455 6.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 4.668 1.14 5.668 1.23 ;
      RECT 5.578 0.891 5.668 1.23 ;
      RECT 5.168 0.875 5.258 1.23 ;
      RECT 4.668 0.53 4.758 1.23 ;
      RECT 5.624 0.846 5.714 0.929 ;
      RECT 5.624 0.846 5.76 0.883 ;
      RECT 5.668 0.801 5.777 0.852 ;
      RECT 5.668 0.801 5.815 0.824 ;
      RECT 5.777 0.715 6.381 0.805 ;
      RECT 5.714 0.755 6.381 0.805 ;
      RECT 5.76 0.723 5.777 0.852 ;
      RECT 4.668 0.53 4.982 0.62 ;
      RECT 4.892 0.35 4.982 0.62 ;
      RECT 4.892 0.35 5.032 0.44 ;
      RECT 5.398 0.275 5.488 1.05 ;
      RECT 5.398 0.275 5.593 0.365 ;
      RECT 0.312 1.06 1.992 1.15 ;
      RECT 0.312 0.25 0.402 1.15 ;
      RECT 4.038 0.25 4.374 0.34 ;
      RECT 2.596 0.25 2.819 0.34 ;
      RECT 0.312 0.25 1.989 0.34 ;
      RECT 4.492 0.17 5.208 0.26 ;
      RECT 2.937 0.17 3.92 0.26 ;
      RECT 2.107 0.17 2.478 0.26 ;
      RECT 5.254 0.17 5.298 0.591 ;
      RECT 5.208 0.17 5.254 0.636 ;
      RECT 5.192 0.534 5.208 0.667 ;
      RECT 5.146 0.565 5.192 0.698 ;
      RECT 5.1 0.611 5.146 0.744 ;
      RECT 5.054 0.657 5.1 0.79 ;
      RECT 5.008 0.703 5.054 0.836 ;
      RECT 4.964 0.748 5.008 0.995 ;
      RECT 4.918 0.793 4.964 0.995 ;
      RECT 4.454 0.17 4.492 0.279 ;
      RECT 4.412 0.191 4.454 0.319 ;
      RECT 4.374 0.231 4.412 0.34 ;
      RECT 4 0.231 4.038 0.34 ;
      RECT 3.958 0.191 4 0.319 ;
      RECT 3.92 0.17 3.958 0.279 ;
      RECT 2.899 0.17 2.937 0.279 ;
      RECT 2.857 0.191 2.899 0.319 ;
      RECT 2.819 0.231 2.857 0.34 ;
      RECT 2.558 0.231 2.596 0.34 ;
      RECT 2.516 0.191 2.558 0.319 ;
      RECT 2.478 0.17 2.516 0.279 ;
      RECT 2.069 0.17 2.107 0.279 ;
      RECT 2.027 0.191 2.069 0.319 ;
      RECT 1.989 0.231 2.027 0.34 ;
      RECT 3.646 1.095 4.051 1.185 ;
      RECT 3.961 0.43 4.051 1.185 ;
      RECT 4.373 0.92 4.573 1.01 ;
      RECT 4.483 0.376 4.573 1.01 ;
      RECT 4.529 0.351 4.573 1.01 ;
      RECT 3.952 0.43 4.051 0.563 ;
      RECT 3.92 0.414 3.952 0.542 ;
      RECT 3.92 0.43 4.573 0.52 ;
      RECT 4.452 0.414 4.573 0.52 ;
      RECT 3.874 0.375 3.92 0.503 ;
      RECT 3.836 0.43 4.573 0.461 ;
      RECT 3.196 0.352 3.874 0.442 ;
      RECT 4.532 0.35 4.782 0.44 ;
      RECT 2.301 0.88 3.376 0.97 ;
      RECT 2.292 0.88 3.376 0.966 ;
      RECT 2.246 0.359 2.336 0.938 ;
      RECT 2.246 0.878 2.339 0.938 ;
      RECT 1.807 0.43 1.897 0.755 ;
      RECT 0.492 0.43 0.582 0.705 ;
      RECT 0.492 0.43 2.336 0.52 ;
      RECT 2.246 0.359 2.441 0.449 ;
  END
END MUX4X6H7R

MACRO MUXI2X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUXI2X0P5H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.92 1.035 2.01 1.48 ;
        RECT 0.325 1.24 0.465 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.92 -0.08 2.01 0.405 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.38 0.61 0.58 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.965 0.625 2.145 0.775 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END B
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.85 0.705 1.47 0.795 ;
        RECT 1.38 0.655 1.47 0.795 ;
        RECT 0.49 1.055 0.94 1.145 ;
        RECT 0.85 0.705 0.94 1.145 ;
        RECT 0.49 0.835 0.58 1.145 ;
        RECT 0.225 0.835 0.58 0.925 ;
      LAYER MET2 ;
        RECT 0.65 0.84 0.75 1.22 ;
      LAYER VIA1 ;
        RECT 0.655 1.055 0.745 1.145 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.03 0.885 1.65 0.975 ;
        RECT 1.56 0.455 1.65 0.975 ;
        RECT 1.28 0.455 1.65 0.545 ;
        RECT 1.28 0.28 1.37 0.545 ;
        RECT 1.03 0.885 1.12 1.12 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.255 1.075 1.83 1.165 ;
      RECT 1.74 0.275 1.83 1.165 ;
      RECT 1.53 0.275 1.83 0.365 ;
      RECT 0.67 0.515 0.76 0.955 ;
      RECT 0.67 0.515 1.03 0.605 ;
      RECT 0.94 0.325 1.03 0.605 ;
      RECT 0.045 1.02 0.185 1.11 ;
      RECT 0.045 0.23 0.135 1.11 ;
      RECT 0.045 0.42 0.493 0.51 ;
      RECT 0.045 0.42 0.539 0.487 ;
      RECT 0.455 0.401 0.585 0.441 ;
      RECT 0.493 0.359 0.585 0.441 ;
      RECT 0.539 0.313 0.631 0.395 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.585 0.267 0.677 0.349 ;
      RECT 0.631 0.221 0.743 0.279 ;
      RECT 0.677 0.184 0.705 0.312 ;
      RECT 0.705 0.17 0.876 0.26 ;
  END
END MUXI2X0P5H7R

MACRO MUXI2X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUXI2X0P7H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.92 1.035 2.01 1.48 ;
        RECT 0.325 1.24 0.465 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.92 -0.08 2.01 0.405 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.38 0.61 0.58 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.965 0.625 2.145 0.775 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END B
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.85 0.705 1.47 0.795 ;
        RECT 1.38 0.655 1.47 0.795 ;
        RECT 0.49 1.055 0.94 1.145 ;
        RECT 0.85 0.705 0.94 1.145 ;
        RECT 0.49 0.835 0.58 1.145 ;
        RECT 0.225 0.835 0.58 0.925 ;
      LAYER MET2 ;
        RECT 0.65 0.84 0.75 1.22 ;
      LAYER VIA1 ;
        RECT 0.655 1.055 0.745 1.145 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.03 0.885 1.65 0.975 ;
        RECT 1.56 0.455 1.65 0.975 ;
        RECT 1.28 0.455 1.65 0.545 ;
        RECT 1.28 0.304 1.37 0.545 ;
        RECT 1.03 0.885 1.12 1.088 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.255 1.065 1.83 1.155 ;
      RECT 1.74 0.353 1.83 1.155 ;
      RECT 1.73 0.28 1.74 0.408 ;
      RECT 1.692 0.353 1.83 0.384 ;
      RECT 1.53 0.275 1.73 0.365 ;
      RECT 1.53 0.308 1.786 0.365 ;
      RECT 0.67 0.515 0.76 0.955 ;
      RECT 0.67 0.515 1.03 0.605 ;
      RECT 0.94 0.325 1.03 0.605 ;
      RECT 0.045 1.02 0.185 1.11 ;
      RECT 0.045 0.23 0.135 1.11 ;
      RECT 0.045 0.42 0.493 0.51 ;
      RECT 0.045 0.42 0.539 0.487 ;
      RECT 0.455 0.401 0.585 0.441 ;
      RECT 0.493 0.359 0.585 0.441 ;
      RECT 0.539 0.313 0.631 0.395 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.585 0.267 0.677 0.349 ;
      RECT 0.631 0.221 0.743 0.279 ;
      RECT 0.677 0.184 0.705 0.312 ;
      RECT 0.705 0.17 0.876 0.26 ;
  END
END MUXI2X0P7H7R

MACRO MUXI2X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUXI2X1H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.92 1.035 2.01 1.48 ;
        RECT 0.325 1.24 0.465 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.908 -0.08 1.998 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.38 0.61 0.58 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.965 0.625 2.145 0.775 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END B
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.85 0.705 1.47 0.795 ;
        RECT 1.38 0.655 1.47 0.795 ;
        RECT 0.49 1.055 0.94 1.145 ;
        RECT 0.85 0.705 0.94 1.145 ;
        RECT 0.49 0.835 0.58 1.145 ;
        RECT 0.225 0.835 0.58 0.925 ;
      LAYER MET2 ;
        RECT 0.65 0.84 0.75 1.22 ;
      LAYER VIA1 ;
        RECT 0.655 1.055 0.745 1.145 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.03 0.885 1.65 0.975 ;
        RECT 1.56 0.455 1.65 0.975 ;
        RECT 1.28 0.455 1.65 0.545 ;
        RECT 1.28 0.28 1.37 0.545 ;
        RECT 1.03 0.885 1.12 1.04 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.244 1.075 1.83 1.165 ;
      RECT 1.74 0.353 1.83 1.165 ;
      RECT 1.73 0.28 1.74 0.408 ;
      RECT 1.692 0.353 1.83 0.384 ;
      RECT 1.505 0.275 1.73 0.365 ;
      RECT 1.505 0.308 1.786 0.365 ;
      RECT 0.67 0.515 0.76 0.955 ;
      RECT 0.67 0.515 1.03 0.605 ;
      RECT 0.94 0.325 1.03 0.605 ;
      RECT 0.045 1.02 0.185 1.11 ;
      RECT 0.045 0.23 0.135 1.11 ;
      RECT 0.045 0.42 0.493 0.51 ;
      RECT 0.045 0.42 0.539 0.487 ;
      RECT 0.455 0.401 0.585 0.441 ;
      RECT 0.493 0.359 0.585 0.441 ;
      RECT 0.539 0.313 0.631 0.395 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.585 0.267 0.677 0.349 ;
      RECT 0.631 0.221 0.743 0.279 ;
      RECT 0.677 0.184 0.705 0.312 ;
      RECT 0.705 0.17 0.876 0.26 ;
  END
END MUXI2X1H7R

MACRO MUXI2X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUXI2X1P4H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.946 1.035 2.036 1.48 ;
        RECT 0.322 1.235 0.465 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.908 -0.08 1.998 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.38 0.61 0.58 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.965 0.625 2.145 0.775 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END B
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.85 0.705 1.47 0.795 ;
        RECT 1.38 0.655 1.47 0.795 ;
        RECT 0.455 1.055 0.94 1.145 ;
        RECT 0.85 0.705 0.94 1.145 ;
        RECT 0.455 0.835 0.545 1.145 ;
        RECT 0.225 0.835 0.545 0.925 ;
      LAYER MET2 ;
        RECT 0.65 0.84 0.75 1.22 ;
      LAYER VIA1 ;
        RECT 0.655 1.055 0.745 1.145 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.03 0.885 1.65 0.975 ;
        RECT 1.56 0.455 1.65 0.975 ;
        RECT 1.28 0.455 1.65 0.545 ;
        RECT 1.28 0.28 1.37 0.545 ;
        RECT 1.03 0.885 1.12 1.03 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.244 1.075 1.83 1.165 ;
      RECT 1.74 0.353 1.83 1.165 ;
      RECT 1.73 0.28 1.74 0.408 ;
      RECT 1.692 0.353 1.83 0.384 ;
      RECT 1.505 0.275 1.73 0.365 ;
      RECT 1.505 0.308 1.786 0.365 ;
      RECT 0.67 0.515 0.76 0.965 ;
      RECT 0.67 0.515 1.03 0.605 ;
      RECT 0.94 0.325 1.03 0.605 ;
      RECT 0.045 1.02 0.185 1.11 ;
      RECT 0.045 0.23 0.135 1.11 ;
      RECT 0.045 0.43 0.483 0.52 ;
      RECT 0.045 0.43 0.529 0.497 ;
      RECT 0.445 0.411 0.575 0.451 ;
      RECT 0.483 0.369 0.575 0.451 ;
      RECT 0.529 0.323 0.621 0.405 ;
      RECT 0.575 0.277 0.667 0.359 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.621 0.231 0.743 0.279 ;
      RECT 0.667 0.189 0.705 0.317 ;
      RECT 0.705 0.17 0.876 0.26 ;
  END
END MUXI2X1P4H7R

MACRO MUXI2X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUXI2X2H7R 0 0 ;
  SIZE 3.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.2 1.48 ;
        RECT 2.945 1.015 3.035 1.48 ;
        RECT 2.425 1.15 2.515 1.48 ;
        RECT 0.31 1.155 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.2 0.08 ;
        RECT 2.94 -0.08 3.03 0.45 ;
        RECT 2.41 -0.08 2.5 0.455 ;
        RECT 0.31 -0.08 0.45 0.245 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.63 0.54 0.77 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.455 0.615 2.62 0.78 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END B
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1 0.77 1.64 0.86 ;
        RECT 1.455 0.615 1.64 0.86 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.93 0.17 2.02 0.35 ;
        RECT 1.35 1.14 1.98 1.23 ;
        RECT 1.32 0.17 2.02 0.26 ;
        RECT 0.805 0.35 1.46 0.44 ;
        RECT 1.32 0.17 1.46 0.44 ;
        RECT 1.35 0.96 1.44 1.23 ;
        RECT 0.805 0.96 1.44 1.05 ;
        RECT 0.805 0.35 0.945 0.575 ;
        RECT 0.805 0.35 0.9 1.05 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.66 0.96 2.805 1.095 ;
      RECT 2.715 0.335 2.805 1.095 ;
      RECT 1.575 0.96 2.805 1.05 ;
      RECT 1.75 0.35 1.84 1.05 ;
      RECT 1.59 0.35 1.84 0.44 ;
      RECT 2.635 0.335 2.805 0.425 ;
      RECT 2.085 0.58 2.25 0.87 ;
      RECT 2.16 0.31 2.25 0.87 ;
      RECT 1.97 0.58 2.25 0.67 ;
      RECT 0.605 1.14 1.235 1.23 ;
      RECT 0.605 0.95 0.695 1.23 ;
      RECT 0.045 0.95 0.695 1.065 ;
      RECT 0.045 0.335 0.135 1.065 ;
      RECT 0.045 0.335 0.69 0.45 ;
      RECT 0.6 0.17 0.69 0.45 ;
      RECT 0.6 0.17 1.23 0.26 ;
  END
END MUXI2X2H7R

MACRO MUXI2X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUXI2X3H7R 0 0 ;
  SIZE 3.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.2 1.48 ;
        RECT 2.945 1.035 3.035 1.48 ;
        RECT 2.425 1.15 2.515 1.48 ;
        RECT 0.31 1.07 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.2 0.08 ;
        RECT 2.94 -0.08 3.03 0.375 ;
        RECT 2.41 -0.08 2.5 0.385 ;
        RECT 0.31 -0.08 0.45 0.335 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.63 0.525 0.77 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.455 0.615 2.62 0.78 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END B
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.62 1.62 0.71 ;
        RECT 1.53 0.57 1.62 0.71 ;
        RECT 1.055 0.62 1.145 0.87 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.915 0.17 2.005 0.39 ;
        RECT 1.35 1.14 1.98 1.23 ;
        RECT 1.35 0.17 2.005 0.26 ;
        RECT 1.35 0.96 1.44 1.23 ;
        RECT 0.855 0.44 1.44 0.53 ;
        RECT 1.35 0.17 1.44 0.53 ;
        RECT 0.855 0.96 1.44 1.05 ;
        RECT 0.815 0.35 0.955 0.44 ;
        RECT 0.855 0.35 0.945 1.05 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.575 0.96 2.805 1.05 ;
      RECT 2.715 0.35 2.805 1.05 ;
      RECT 1.735 0.35 1.825 1.05 ;
      RECT 2.635 0.35 2.805 0.44 ;
      RECT 1.59 0.35 1.825 0.44 ;
      RECT 2.105 0.58 2.25 0.87 ;
      RECT 2.16 0.31 2.25 0.87 ;
      RECT 1.97 0.58 2.25 0.67 ;
      RECT 0.59 1.14 1.235 1.23 ;
      RECT 0.59 0.89 0.68 1.23 ;
      RECT 0.045 0.89 0.185 1.01 ;
      RECT 0.045 0.89 0.68 0.98 ;
      RECT 0.045 0.335 0.135 1.01 ;
      RECT 0.045 0.425 0.675 0.515 ;
      RECT 0.585 0.17 0.675 0.515 ;
      RECT 0.045 0.335 0.185 0.515 ;
      RECT 1.095 0.17 1.235 0.35 ;
      RECT 0.585 0.17 1.235 0.26 ;
  END
END MUXI2X3H7R

MACRO MUXI2X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUXI2X4H7R 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.8 1.48 ;
        RECT 3.291 1.105 3.431 1.48 ;
        RECT 2.761 1.225 2.901 1.48 ;
        RECT 0.31 1.075 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.8 0.08 ;
        RECT 3.255 -0.08 3.345 0.245 ;
        RECT 2.74 -0.08 2.83 0.385 ;
        RECT 0.575 -0.08 0.715 0.175 ;
        RECT 0.045 -0.08 0.185 0.175 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.645 0.79 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.895 0.655 3.435 0.745 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END B
  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.545 1.915 0.635 ;
        RECT 1.285 0.71 1.545 0.8 ;
        RECT 1.455 0.545 1.545 0.8 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.2 0.17 2.29 0.39 ;
        RECT 1.645 1.095 2.26 1.185 ;
        RECT 1.69 0.17 2.29 0.26 ;
        RECT 1.055 0.35 1.78 0.44 ;
        RECT 1.69 0.17 1.78 0.44 ;
        RECT 1.645 0.895 1.735 1.185 ;
        RECT 1.055 0.895 1.735 0.985 ;
        RECT 1.055 0.35 1.145 0.985 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.426 1.04 3.116 1.13 ;
      RECT 3.026 0.925 3.116 1.13 ;
      RECT 2.411 0.994 2.426 1.123 ;
      RECT 2.365 0.964 2.411 1.092 ;
      RECT 2.319 0.918 2.365 1.046 ;
      RECT 2.319 1.021 2.464 1.046 ;
      RECT 3.026 0.925 3.671 1.015 ;
      RECT 3.581 0.335 3.671 1.015 ;
      RECT 2.281 0.895 2.319 1.004 ;
      RECT 1.87 0.895 2.319 0.985 ;
      RECT 2.005 0.35 2.095 0.985 ;
      RECT 1.925 0.35 2.095 0.44 ;
      RECT 2.965 0.335 3.671 0.425 ;
      RECT 2.501 0.31 2.591 0.949 ;
      RECT 2.3 0.58 2.591 0.67 ;
      RECT 2.49 0.31 2.591 0.67 ;
      RECT 0.58 1.075 1.495 1.165 ;
      RECT 0.58 0.875 0.92 1.165 ;
      RECT 0.045 0.875 0.92 0.965 ;
      RECT 0.045 0.265 0.135 0.965 ;
      RECT 0.045 0.265 0.955 0.355 ;
      RECT 0.865 0.17 0.955 0.355 ;
      RECT 0.865 0.17 1.54 0.26 ;
  END
END MUXI2X4H7R

MACRO NAND2BX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BX0P5H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.81 1.125 0.95 1.48 ;
        RECT 0.295 0.975 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.295 -0.08 0.435 0.32 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.43 0.575 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.65 0.41 0.76 0.66 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.545 0.945 0.945 1.035 ;
        RECT 0.855 0.23 0.945 1.035 ;
        RECT 0.765 0.23 0.945 0.32 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.205 0.16 1.075 ;
      RECT 0.07 0.72 0.545 0.81 ;
  END
END NAND2BX0P5H7R

MACRO NAND2BX0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BX0P7H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.815 1.095 0.955 1.48 ;
        RECT 0.32 0.95 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.43 0.58 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.615 0.425 0.765 0.605 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 0.915 0.945 1.005 ;
        RECT 0.855 0.245 0.945 1.005 ;
        RECT 0.77 0.245 0.945 0.335 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.055 0.205 0.16 1.035 ;
      RECT 0.055 0.703 0.575 0.793 ;
  END
END NAND2BX0P7H7R

MACRO NAND2BX12H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BX12H7R 0 0 ;
  SIZE 4.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.4 1.48 ;
        RECT 3.765 1.07 3.855 1.48 ;
        RECT 3.265 1.07 3.355 1.48 ;
        RECT 2.765 1.07 2.855 1.48 ;
        RECT 2.265 1.07 2.355 1.48 ;
        RECT 1.765 1.07 1.855 1.48 ;
        RECT 1.265 1.07 1.355 1.48 ;
        RECT 0.535 1.07 0.625 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.4 0.08 ;
        RECT 2.24 -0.08 2.38 0.305 ;
        RECT 1.74 -0.08 1.88 0.305 ;
        RECT 1.24 -0.08 1.38 0.305 ;
        RECT 0.51 -0.08 0.65 0.305 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.355 0.655 0.695 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.725 0.655 3.865 0.745 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.015 0.855 4.145 0.945 ;
        RECT 4.055 0.395 4.145 0.945 ;
        RECT 4.015 0.855 4.105 1.195 ;
        RECT 2.74 0.395 4.145 0.485 ;
        RECT 3.515 0.855 3.605 1.2 ;
        RECT 3.015 0.855 3.105 1.2 ;
        RECT 2.515 0.855 2.605 1.2 ;
        RECT 2.015 0.855 2.105 1.2 ;
        RECT 1.515 0.855 1.605 1.2 ;
        RECT 1.015 0.855 1.105 1.195 ;
      LAYER MET2 ;
        RECT 4.05 0.23 4.15 0.76 ;
      LAYER VIA1 ;
        RECT 4.055 0.455 4.145 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.015 0.395 2.605 0.485 ;
      RECT 2.515 0.215 2.605 0.485 ;
      RECT 1.015 0.345 1.105 0.485 ;
      RECT 2.515 0.215 4.13 0.305 ;
      RECT 0.26 0.875 0.875 0.965 ;
      RECT 0.785 0.355 0.875 0.965 ;
      RECT 0.785 0.655 2.34 0.745 ;
      RECT 0.285 0.395 0.875 0.485 ;
      RECT 0.285 0.32 0.375 0.485 ;
  END
END NAND2BX12H7R

MACRO NAND2BX16H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BX16H7R 0 0 ;
  SIZE 7 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7 1.48 ;
        RECT 6.28 1.07 6.37 1.48 ;
        RECT 5.78 1.055 5.87 1.48 ;
        RECT 5.28 1.07 5.37 1.48 ;
        RECT 4.78 1.07 4.87 1.48 ;
        RECT 4.28 1.07 4.37 1.48 ;
        RECT 3.78 1.07 3.87 1.48 ;
        RECT 3.28 1.07 3.37 1.48 ;
        RECT 2.78 1.07 2.87 1.48 ;
        RECT 2.035 1.07 2.125 1.48 ;
        RECT 1.535 1.07 1.625 1.48 ;
        RECT 1.035 1.07 1.125 1.48 ;
        RECT 0.535 1.07 0.625 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7 0.08 ;
        RECT 4.255 -0.08 4.395 0.305 ;
        RECT 3.755 -0.08 3.895 0.305 ;
        RECT 3.255 -0.08 3.395 0.305 ;
        RECT 2.755 -0.08 2.895 0.305 ;
        RECT 2.01 -0.08 2.15 0.305 ;
        RECT 1.51 -0.08 1.65 0.305 ;
        RECT 1.01 -0.08 1.15 0.305 ;
        RECT 0.51 -0.08 0.65 0.305 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.46 0.655 2.215 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.7 0.655 6.44 0.745 ;
      LAYER MET2 ;
        RECT 5.85 0.43 5.95 0.96 ;
      LAYER VIA1 ;
        RECT 5.855 0.655 5.945 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.53 0.395 6.62 1.165 ;
        RECT 2.53 0.855 6.62 0.945 ;
        RECT 4.745 0.395 6.62 0.485 ;
        RECT 6.03 0.855 6.12 1.2 ;
        RECT 5.53 0.855 5.62 1.2 ;
        RECT 5.03 0.855 5.12 1.2 ;
        RECT 4.53 0.855 4.62 1.17 ;
        RECT 4.03 0.855 4.12 1.17 ;
        RECT 3.53 0.855 3.62 1.17 ;
        RECT 3.03 0.855 3.12 1.17 ;
        RECT 2.53 0.855 2.62 1.195 ;
      LAYER MET2 ;
        RECT 6.45 0.625 6.55 1.16 ;
      LAYER VIA1 ;
        RECT 6.455 0.855 6.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.53 0.395 4.62 0.485 ;
      RECT 4.53 0.215 4.62 0.485 ;
      RECT 2.53 0.345 2.62 0.485 ;
      RECT 4.53 0.215 6.645 0.305 ;
      RECT 0.26 0.885 2.4 0.975 ;
      RECT 2.31 0.395 2.4 0.975 ;
      RECT 2.31 0.625 4.44 0.715 ;
      RECT 0.285 0.395 2.4 0.485 ;
      RECT 0.285 0.32 0.375 0.485 ;
  END
END NAND2BX16H7R

MACRO NAND2BX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BX1H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.815 1.145 0.955 1.48 ;
        RECT 0.295 0.96 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.325 -0.08 0.465 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.38 0.635 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.5 0.775 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.545 0.96 0.955 1.05 ;
        RECT 0.865 0.225 0.955 1.05 ;
        RECT 0.84 0.225 0.955 0.375 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.56 ;
      LAYER VIA1 ;
        RECT 0.855 0.255 0.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.285 0.16 1.09 ;
      RECT 0.07 0.73 0.555 0.87 ;
  END
END NAND2BX1H7R

MACRO NAND2BX1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BX1P4H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.8 1.095 0.94 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.41 0.595 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.51 0.775 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 0.915 0.955 1.005 ;
        RECT 0.865 0.225 0.955 1.005 ;
        RECT 0.84 0.225 0.955 0.375 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.56 ;
      LAYER VIA1 ;
        RECT 0.855 0.255 0.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.205 0.16 1.155 ;
      RECT 0.07 0.725 0.545 0.815 ;
  END
END NAND2BX1P4H7R

MACRO NAND2BX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BX2H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.34 1.2 1.48 1.48 ;
        RECT 0.81 1.2 0.95 1.48 ;
        RECT 0.295 1.075 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.34 -0.08 1.48 0.31 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.385 0.625 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.615 1.035 0.705 ;
        RECT 0.655 0.425 0.745 0.705 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.545 1.005 1.545 1.095 ;
        RECT 1.455 0.435 1.545 1.095 ;
        RECT 0.835 0.435 1.545 0.525 ;
        RECT 0.835 0.215 0.925 0.525 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.205 0.16 1.135 ;
      RECT 0.07 0.8 1.365 0.89 ;
  END
END NAND2BX2H7R

MACRO NAND2BX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BX3H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.325 1.075 1.465 1.48 ;
        RECT 0.81 1.075 0.95 1.48 ;
        RECT 0.32 1.05 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.39 -0.08 1.53 0.185 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.385 0.625 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.725 0.455 1.065 0.58 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.57 0.895 1.545 0.985 ;
        RECT 1.455 0.275 1.545 0.985 ;
        RECT 0.825 0.275 1.545 0.365 ;
        RECT 1.1 0.895 1.19 1.04 ;
        RECT 0.57 0.895 0.66 1.04 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.205 0.16 1.135 ;
      RECT 0.07 0.715 1.315 0.805 ;
  END
END NAND2BX3H7R

MACRO NAND2BX4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BX4H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 2.375 1.075 2.515 1.48 ;
        RECT 1.875 1.075 2.015 1.48 ;
        RECT 1.345 1.075 1.485 1.48 ;
        RECT 0.845 1.075 0.985 1.48 ;
        RECT 0.33 0.9 0.47 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 2.39 -0.08 2.53 0.175 ;
        RECT 1.36 -0.08 1.5 0.175 ;
        RECT 0.325 -0.08 0.465 0.325 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.455 0.575 0.605 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.745 0.495 2.115 0.585 ;
        RECT 1.425 0.455 1.575 0.585 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.595 0.895 2.545 0.985 ;
        RECT 2.455 0.265 2.545 0.985 ;
        RECT 0.845 0.265 2.545 0.355 ;
        RECT 2.125 0.895 2.265 1.095 ;
        RECT 1.625 0.895 1.765 1.095 ;
        RECT 1.095 0.895 1.235 1.095 ;
        RECT 0.595 0.895 0.735 1.095 ;
      LAYER MET2 ;
        RECT 2.45 0.625 2.55 1.16 ;
      LAYER VIA1 ;
        RECT 2.455 0.855 2.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.265 0.16 1.215 ;
      RECT 0.07 0.715 2.365 0.805 ;
  END
END NAND2BX4H7R

MACRO NAND2BX6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BX6H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 2.035 1.055 2.125 1.48 ;
        RECT 1.535 1.07 1.625 1.48 ;
        RECT 1.035 1.07 1.125 1.48 ;
        RECT 0.535 1.07 0.625 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 1.01 -0.08 1.15 0.305 ;
        RECT 0.535 -0.08 0.625 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.425 0.545 0.71 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.425 0.655 1.965 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.785 0.86 2.145 0.95 ;
        RECT 2.055 0.315 2.145 0.95 ;
        RECT 1.51 0.395 2.145 0.485 ;
        RECT 1.785 0.86 1.875 1.2 ;
        RECT 1.285 0.86 1.375 1.2 ;
        RECT 0.785 0.86 0.875 1.2 ;
      LAYER MET2 ;
        RECT 2.05 0.23 2.15 0.76 ;
      LAYER VIA1 ;
        RECT 2.055 0.455 2.145 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.76 0.395 1.375 0.485 ;
      RECT 1.285 0.215 1.375 0.485 ;
      RECT 1.285 0.215 1.9 0.305 ;
      RECT 0.26 0.875 0.375 1.19 ;
      RECT 0.26 0.875 0.549 0.965 ;
      RECT 0.26 0.875 0.595 0.942 ;
      RECT 0.511 0.856 0.641 0.896 ;
      RECT 0.26 0.23 0.355 1.19 ;
      RECT 0.549 0.814 0.641 0.896 ;
      RECT 0.549 0.814 0.687 0.85 ;
      RECT 0.595 0.768 0.69 0.826 ;
      RECT 0.641 0.722 0.736 0.801 ;
      RECT 0.687 0.697 0.69 0.826 ;
      RECT 0.641 0.722 0.769 0.762 ;
      RECT 0.69 0.655 1.23 0.745 ;
      RECT 0.26 0.23 0.4 0.32 ;
  END
END NAND2BX6H7R

MACRO NAND2BX8H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BX8H7R 0 0 ;
  SIZE 3.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.2 1.48 ;
        RECT 2.815 1.055 2.905 1.48 ;
        RECT 2.315 1.07 2.405 1.48 ;
        RECT 1.815 1.07 1.905 1.48 ;
        RECT 1.315 1.07 1.405 1.48 ;
        RECT 0.815 1.055 0.905 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.2 0.08 ;
        RECT 1.54 -0.08 1.68 0.305 ;
        RECT 1.04 -0.08 1.18 0.305 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.195 0.655 0.535 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.97 0.655 2.715 0.745 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.065 0.87 2.945 0.96 ;
        RECT 2.855 0.395 2.945 0.96 ;
        RECT 2.04 0.395 2.945 0.485 ;
        RECT 2.565 0.87 2.655 1.21 ;
        RECT 2.065 0.87 2.155 1.21 ;
        RECT 1.565 0.87 1.655 1.21 ;
        RECT 1.065 0.87 1.155 1.21 ;
      LAYER MET2 ;
        RECT 2.85 0.23 2.95 0.76 ;
      LAYER VIA1 ;
        RECT 2.855 0.455 2.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.815 0.395 1.905 0.485 ;
      RECT 1.815 0.215 1.905 0.485 ;
      RECT 0.815 0.345 0.905 0.485 ;
      RECT 1.815 0.215 2.93 0.305 ;
      RECT 0.07 0.915 0.16 1.06 ;
      RECT 0.07 0.915 0.715 1.005 ;
      RECT 0.625 0.496 0.715 1.005 ;
      RECT 0.625 0.655 1.71 0.745 ;
      RECT 0.617 0.496 0.715 0.535 ;
      RECT 0.571 0.469 0.706 0.508 ;
      RECT 0.57 0.305 0.66 0.485 ;
      RECT 0.07 0.395 0.66 0.485 ;
      RECT 0.07 0.305 0.16 0.485 ;
  END
END NAND2BX8H7R

MACRO NAND2X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X0P5H7R 0 0 ;
  SIZE 0.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.8 1.48 ;
        RECT 0.555 1.075 0.695 1.48 ;
        RECT 0.07 1.05 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.8 0.08 ;
        RECT 0.045 -0.08 0.185 0.32 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.505 0.625 0.745 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.425 0.23 0.685 ;
      LAYER MET2 ;
        RECT 0.05 0.23 0.15 0.76 ;
      LAYER VIA1 ;
        RECT 0.055 0.455 0.145 0.545 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.32 0.23 0.685 0.32 ;
        RECT 0.32 0.23 0.41 1.14 ;
        RECT 0.255 0.825 0.41 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END Y
END NAND2X0P5H7R

MACRO NAND2X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X0P7H7R 0 0 ;
  SIZE 0.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.8 1.48 ;
        RECT 0.57 1.055 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.8 0.08 ;
        RECT 0.045 -0.08 0.185 0.32 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.425 0.23 0.58 ;
      LAYER MET2 ;
        RECT 0.05 0.23 0.15 0.76 ;
      LAYER VIA1 ;
        RECT 0.055 0.455 0.145 0.545 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.5 0.625 0.745 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.32 0.255 0.685 0.345 ;
        RECT 0.32 0.255 0.41 1.108 ;
        RECT 0.255 0.825 0.41 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END Y
END NAND2X0P7H7R

MACRO NAND2X12H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X12H7R 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.8 1.48 ;
        RECT 3.325 1.07 3.415 1.48 ;
        RECT 2.825 1.07 2.915 1.48 ;
        RECT 2.325 1.07 2.415 1.48 ;
        RECT 1.825 1.07 1.915 1.48 ;
        RECT 1.325 1.07 1.415 1.48 ;
        RECT 0.825 1.07 0.915 1.48 ;
        RECT 0.325 1.055 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.8 0.08 ;
        RECT 1.55 -0.08 1.69 0.305 ;
        RECT 1.05 -0.08 1.19 0.305 ;
        RECT 0.55 -0.08 0.69 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.98 0.655 3.12 0.745 ;
      LAYER MET2 ;
        RECT 2.85 0.43 2.95 0.96 ;
      LAYER VIA1 ;
        RECT 2.855 0.655 2.945 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.495 0.655 1.635 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 0.885 3.345 0.975 ;
        RECT 3.255 0.395 3.345 0.975 ;
        RECT 2.05 0.395 3.345 0.485 ;
      LAYER MET2 ;
        RECT 3.25 0.63 3.35 1.16 ;
      LAYER VIA1 ;
        RECT 3.255 0.855 3.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.325 0.395 1.94 0.485 ;
      RECT 1.85 0.215 1.94 0.485 ;
      RECT 0.325 0.345 0.415 0.485 ;
      RECT 1.85 0.215 3.44 0.305 ;
  END
END NAND2X12H7R

MACRO NAND2X16H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X16H7R 0 0 ;
  SIZE 4.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.8 1.48 ;
        RECT 4.325 1.07 4.415 1.48 ;
        RECT 3.825 1.07 3.915 1.48 ;
        RECT 3.325 1.07 3.415 1.48 ;
        RECT 2.825 1.07 2.915 1.48 ;
        RECT 2.325 1.07 2.415 1.48 ;
        RECT 1.825 1.07 1.915 1.48 ;
        RECT 1.325 1.07 1.415 1.48 ;
        RECT 0.825 1.07 0.915 1.48 ;
        RECT 0.325 1.055 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.8 0.08 ;
        RECT 2.05 -0.08 2.19 0.305 ;
        RECT 1.55 -0.08 1.69 0.305 ;
        RECT 1.05 -0.08 1.19 0.305 ;
        RECT 0.55 -0.08 0.69 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.5 0.655 4.24 0.745 ;
      LAYER MET2 ;
        RECT 3.85 0.43 3.95 0.96 ;
      LAYER VIA1 ;
        RECT 3.855 0.655 3.945 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.495 0.655 2.235 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 0.885 4.545 0.975 ;
        RECT 4.455 0.395 4.545 0.975 ;
        RECT 2.55 0.395 4.545 0.485 ;
      LAYER MET2 ;
        RECT 4.45 0.625 4.55 1.16 ;
      LAYER VIA1 ;
        RECT 4.455 0.855 4.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.325 0.395 2.44 0.485 ;
      RECT 2.35 0.215 2.44 0.485 ;
      RECT 0.325 0.345 0.415 0.485 ;
      RECT 2.35 0.215 4.44 0.305 ;
  END
END NAND2X16H7R

MACRO NAND2X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X1H7R 0 0 ;
  SIZE 0.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.8 1.48 ;
        RECT 0.555 1.075 0.695 1.48 ;
        RECT 0.045 1.075 0.185 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.8 0.08 ;
        RECT 0.045 -0.08 0.185 0.325 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.425 0.23 0.59 ;
      LAYER MET2 ;
        RECT 0.05 0.23 0.15 0.76 ;
      LAYER VIA1 ;
        RECT 0.055 0.455 0.145 0.545 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.5 0.625 0.745 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.32 0.285 0.685 0.375 ;
        RECT 0.32 0.285 0.41 1.09 ;
        RECT 0.255 0.825 0.41 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END Y
END NAND2X1H7R

MACRO NAND2X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X1P4H7R 0 0 ;
  SIZE 0.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.8 1.48 ;
        RECT 0.57 1.055 0.66 1.48 ;
        RECT 0.045 1.08 0.185 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.8 0.08 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.825 0.23 0.975 ;
        RECT 0.14 0.7 0.23 0.975 ;
      LAYER MET2 ;
        RECT 0.05 0.625 0.15 1.16 ;
      LAYER VIA1 ;
        RECT 0.055 0.855 0.145 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.5 0.625 0.745 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.32 0.326 0.685 0.416 ;
        RECT 0.32 0.326 0.41 1.016 ;
        RECT 0.255 0.425 0.41 0.575 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END Y
END NAND2X1P4H7R

MACRO NAND2X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X2H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.165 1.055 1.255 1.48 ;
        RECT 0.63 1.095 0.77 1.48 ;
        RECT 0.105 1.055 0.195 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.345 -0.08 0.485 0.225 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.545 0.765 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.815 0.68 1.345 0.82 ;
        RECT 1.255 0.625 1.345 0.82 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.635 0.5 1.03 0.59 ;
        RECT 0.89 0.35 1.03 0.59 ;
        RECT 0.915 0.915 1.005 1.14 ;
        RECT 0.355 0.915 1.005 1.005 ;
        RECT 0.355 0.855 0.725 1.005 ;
        RECT 0.635 0.5 0.725 1.005 ;
        RECT 0.355 0.855 0.445 1.145 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.165 0.17 1.255 0.45 ;
      RECT 0.08 0.32 0.755 0.41 ;
      RECT 0.665 0.17 0.755 0.41 ;
      RECT 0.665 0.17 1.255 0.26 ;
  END
END NAND2X2H7R

MACRO NAND2X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X3H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.165 1.055 1.255 1.48 ;
        RECT 0.63 1.095 0.77 1.48 ;
        RECT 0.105 1.055 0.195 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.345 -0.08 0.485 0.175 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.655 0.565 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.835 0.655 1.175 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.445 1.03 0.535 ;
        RECT 0.89 0.35 1.03 0.535 ;
        RECT 0.915 0.905 1.005 1.045 ;
        RECT 0.355 0.905 1.005 0.995 ;
        RECT 0.655 0.445 0.745 0.995 ;
        RECT 0.355 0.905 0.445 1.045 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.165 0.17 1.255 0.375 ;
      RECT 0.08 0.265 0.755 0.355 ;
      RECT 0.64 0.17 0.755 0.355 ;
      RECT 0.64 0.17 1.255 0.26 ;
  END
END NAND2X3H7R

MACRO NAND2X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X4H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 2.215 1.08 2.355 1.48 ;
        RECT 1.715 1.095 1.855 1.48 ;
        RECT 1.065 1.095 1.205 1.48 ;
        RECT 0.545 1.095 0.685 1.48 ;
        RECT 0.045 1.08 0.185 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 0.795 -0.08 0.935 0.41 ;
        RECT 0.295 -0.08 0.435 0.41 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.69 0.965 0.78 ;
        RECT 0.055 0.69 0.145 0.975 ;
      LAYER MET2 ;
        RECT 0.05 0.625 0.15 1.16 ;
      LAYER VIA1 ;
        RECT 0.055 0.855 0.145 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.435 0.69 2.345 0.78 ;
        RECT 2.255 0.625 2.345 0.78 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.965 0.915 2.105 1.115 ;
        RECT 1.255 0.5 2.105 0.59 ;
        RECT 1.965 0.35 2.105 0.59 ;
        RECT 0.295 0.915 2.105 1.005 ;
        RECT 1.465 0.915 1.605 1.115 ;
        RECT 1.465 0.35 1.605 0.59 ;
        RECT 1.255 0.5 1.345 1.005 ;
        RECT 0.795 0.915 0.935 1.115 ;
        RECT 0.295 0.915 0.435 1.12 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.5 1.16 0.59 ;
      RECT 1.07 0.17 1.16 0.59 ;
      RECT 0.545 0.35 0.685 0.59 ;
      RECT 0.045 0.335 0.185 0.59 ;
      RECT 2.215 0.17 2.355 0.425 ;
      RECT 1.715 0.17 1.855 0.41 ;
      RECT 1.07 0.17 2.355 0.26 ;
  END
END NAND2X4H7R

MACRO NAND2X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X6H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.785 1.07 1.875 1.48 ;
        RECT 1.285 1.07 1.375 1.48 ;
        RECT 0.785 1.07 0.875 1.48 ;
        RECT 0.285 1.055 0.375 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 0.76 -0.08 0.9 0.305 ;
        RECT 0.285 -0.08 0.375 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.175 0.655 1.715 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.43 0.655 0.97 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.51 0.885 1.945 0.975 ;
        RECT 1.855 0.395 1.945 0.975 ;
        RECT 1.785 0.31 1.875 0.485 ;
        RECT 1.26 0.395 1.945 0.485 ;
      LAYER MET2 ;
        RECT 1.85 0.625 1.95 1.16 ;
      LAYER VIA1 ;
        RECT 1.855 0.855 1.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.51 0.395 1.15 0.485 ;
      RECT 1.06 0.215 1.15 0.485 ;
      RECT 1.06 0.215 1.65 0.305 ;
  END
END NAND2X6H7R

MACRO NAND2X8H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X8H7R 0 0 ;
  SIZE 2.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.8 1.48 ;
        RECT 2.325 1.07 2.415 1.48 ;
        RECT 1.825 1.07 1.915 1.48 ;
        RECT 1.325 1.07 1.415 1.48 ;
        RECT 0.825 1.07 0.915 1.48 ;
        RECT 0.325 1.055 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.8 0.08 ;
        RECT 1.05 -0.08 1.19 0.305 ;
        RECT 0.55 -0.08 0.69 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.5 0.655 2.24 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.495 0.655 1.235 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 0.885 2.545 0.975 ;
        RECT 2.455 0.395 2.545 0.975 ;
        RECT 1.55 0.395 2.545 0.485 ;
      LAYER MET2 ;
        RECT 2.45 0.625 2.55 1.16 ;
      LAYER VIA1 ;
        RECT 2.455 0.855 2.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.325 0.395 1.44 0.485 ;
      RECT 1.35 0.215 1.44 0.485 ;
      RECT 0.325 0.315 0.415 0.485 ;
      RECT 1.35 0.215 2.44 0.305 ;
  END
END NAND2X8H7R

MACRO NAND3BBX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BBX0P5H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.555 1.055 1.645 1.48 ;
        RECT 0.795 1.095 0.935 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.56 -0.08 1.65 0.345 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.385 0.625 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.565 0.625 1.745 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.575 0.99 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.91 1.175 1.175 ;
        RECT 1.085 0.35 1.175 1.175 ;
        RECT 1.035 0.35 1.175 0.44 ;
        RECT 0.57 0.91 1.175 1 ;
        RECT 0.57 0.91 0.66 1.14 ;
      LAYER MET2 ;
        RECT 1.05 0.84 1.15 1.22 ;
      LAYER VIA1 ;
        RECT 1.055 1.055 1.145 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.305 0.17 1.395 1.155 ;
      RECT 0.67 0.17 0.76 0.555 ;
      RECT 0.67 0.17 1.395 0.26 ;
      RECT 0.07 0.205 0.16 1.155 ;
      RECT 0.07 0.73 0.585 0.82 ;
  END
END NAND3BBX0P5H7R

MACRO NAND3BBX0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BBX0P7H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.565 1.055 1.655 1.48 ;
        RECT 0.795 1.095 0.935 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.57 -0.08 1.66 0.345 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.42 0.385 0.62 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.565 0.625 1.745 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.595 0.99 0.795 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.91 1.175 1.175 ;
        RECT 1.085 0.35 1.175 1.175 ;
        RECT 1.035 0.35 1.175 0.44 ;
        RECT 0.57 0.91 1.175 1 ;
        RECT 0.57 0.91 0.66 1.108 ;
      LAYER MET2 ;
        RECT 1.05 0.84 1.15 1.22 ;
      LAYER VIA1 ;
        RECT 1.055 1.055 1.145 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.315 0.17 1.405 1.155 ;
      RECT 0.67 0.17 0.76 0.58 ;
      RECT 0.67 0.17 1.405 0.26 ;
      RECT 0.07 0.205 0.16 1.16 ;
      RECT 0.07 0.73 0.585 0.82 ;
  END
END NAND3BBX0P7H7R

MACRO NAND3BBX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BBX1H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.32 1.07 1.41 1.48 ;
        RECT 0.79 1.095 0.93 1.48 ;
        RECT 0.32 1.055 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.32 -0.08 1.41 0.33 ;
        RECT 0.32 -0.08 0.41 0.345 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.455 0.375 0.635 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.395 0.795 1.545 0.975 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.175 0.655 1.265 0.825 ;
        RECT 1.025 0.655 1.265 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.065 0.915 1.155 1.06 ;
        RECT 0.55 0.915 1.155 1.005 ;
        RECT 0.845 0.825 0.96 1.005 ;
        RECT 0.845 0.683 0.935 1.005 ;
        RECT 0.778 0.638 0.891 0.699 ;
        RECT 0.732 0.604 0.845 0.653 ;
        RECT 0.824 0.683 0.935 0.733 ;
        RECT 0.686 0.571 0.824 0.607 ;
        RECT 0.686 0.525 0.778 0.607 ;
        RECT 0.64 0.479 0.732 0.561 ;
        RECT 0.596 0.433 0.686 0.516 ;
        RECT 0.55 0.915 0.64 1.075 ;
        RECT 0.55 0.26 0.64 0.471 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.545 1.065 1.725 1.155 ;
      RECT 1.635 0.23 1.725 1.155 ;
      RECT 0.935 0.475 1.725 0.565 ;
      RECT 1.545 0.23 1.725 0.32 ;
      RECT 0.045 1.045 0.185 1.135 ;
      RECT 0.045 0.23 0.135 1.135 ;
      RECT 0.045 0.735 0.705 0.825 ;
      RECT 0.045 0.23 0.185 0.32 ;
  END
END NAND3BBX1H7R

MACRO NAND3BBX1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BBX1P4H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.32 1.07 1.41 1.48 ;
        RECT 0.79 1.095 0.93 1.48 ;
        RECT 0.32 1.055 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.32 -0.08 1.41 0.345 ;
        RECT 0.295 -0.08 0.435 0.32 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.415 0.385 0.615 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.715 1.56 0.975 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.215 0.625 1.35 0.825 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.54 0.915 1.18 1.005 ;
        RECT 0.805 0.255 0.895 1.005 ;
        RECT 0.525 0.255 0.895 0.345 ;
      LAYER MET2 ;
        RECT 0.65 0.18 0.75 0.56 ;
      LAYER VIA1 ;
        RECT 0.655 0.255 0.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.545 1.065 1.74 1.155 ;
      RECT 1.65 0.445 1.74 1.155 ;
      RECT 0.99 0.445 1.08 0.655 ;
      RECT 0.99 0.445 1.74 0.535 ;
      RECT 1.57 0.205 1.66 0.535 ;
      RECT 0.07 0.205 0.16 1.155 ;
      RECT 0.07 0.705 0.715 0.795 ;
  END
END NAND3BBX1P4H7R

MACRO NAND3BBX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BBX2H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.32 1.07 1.41 1.48 ;
        RECT 0.815 1.07 0.905 1.48 ;
        RECT 0.32 1.055 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.32 -0.08 1.41 0.33 ;
        RECT 0.32 -0.08 0.41 0.345 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.455 0.405 0.605 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.395 0.615 1.545 0.795 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.655 1.3 0.755 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.525 0.875 1.18 0.965 ;
        RECT 0.775 0.23 0.865 0.965 ;
        RECT 0.525 0.23 0.865 0.345 ;
      LAYER MET2 ;
        RECT 0.65 0.18 0.75 0.56 ;
      LAYER VIA1 ;
        RECT 0.655 0.255 0.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.545 0.885 1.725 0.975 ;
      RECT 1.635 0.23 1.725 0.975 ;
      RECT 0.955 0.42 1.045 0.56 ;
      RECT 0.955 0.42 1.725 0.51 ;
      RECT 1.545 0.23 1.725 0.32 ;
      RECT 0.045 0.695 0.16 0.965 ;
      RECT 0.045 0.695 0.685 0.785 ;
      RECT 0.595 0.615 0.685 0.785 ;
      RECT 0.045 0.23 0.135 0.965 ;
      RECT 0.045 0.23 0.185 0.32 ;
  END
END NAND3BBX2H7R

MACRO NAND3BBX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BBX3H7R 0 0 ;
  SIZE 2.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.8 1.48 ;
        RECT 2.37 1.07 2.46 1.48 ;
        RECT 1.61 1.07 1.7 1.48 ;
        RECT 1.08 1.07 1.17 1.48 ;
        RECT 0.55 1.055 0.64 1.48 ;
        RECT 0.32 1.055 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.8 0.08 ;
        RECT 2.37 -0.08 2.46 0.33 ;
        RECT 1.845 -0.08 1.985 0.305 ;
        RECT 0.32 -0.08 0.41 0.345 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.455 0.405 0.605 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.435 0.775 2.57 0.975 ;
      LAYER MET2 ;
        RECT 2.45 0.625 2.55 1.16 ;
      LAYER VIA1 ;
        RECT 2.455 0.855 2.545 0.945 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.995 0.76 2.335 0.85 ;
        RECT 1.995 0.76 2.175 0.945 ;
      LAYER MET2 ;
        RECT 2.05 0.63 2.15 1.16 ;
      LAYER VIA1 ;
        RECT 2.055 0.855 2.145 0.945 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.79 1.055 2.235 1.145 ;
        RECT 1.79 0.89 1.88 1.145 ;
        RECT 0.8 0.89 1.88 0.98 ;
        RECT 1.305 0.89 1.445 1.02 ;
        RECT 0.885 0.35 0.975 0.98 ;
        RECT 0.8 0.89 0.89 1.045 ;
        RECT 0.79 0.35 0.975 0.44 ;
      LAYER MET2 ;
        RECT 1.85 0.84 1.95 1.22 ;
      LAYER VIA1 ;
        RECT 1.855 1.055 1.945 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.595 1.065 2.75 1.155 ;
      RECT 2.66 0.23 2.75 1.155 ;
      RECT 1.235 0.58 2.75 0.67 ;
      RECT 2.595 0.23 2.75 0.32 ;
      RECT 1.32 0.4 2.21 0.49 ;
      RECT 2.12 0.295 2.21 0.49 ;
      RECT 1.32 0.35 1.46 0.49 ;
      RECT 0.55 0.17 0.64 0.345 ;
      RECT 1.585 0.17 1.725 0.305 ;
      RECT 1.055 0.17 1.195 0.305 ;
      RECT 0.55 0.17 1.725 0.26 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 0.045 0.71 0.79 0.8 ;
      RECT 0.7 0.66 0.79 0.8 ;
      RECT 0.045 0.23 0.185 0.32 ;
  END
END NAND3BBX3H7R

MACRO NAND3BBX4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BBX4H7R 0 0 ;
  SIZE 2.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.8 1.48 ;
        RECT 2.57 1.055 2.66 1.48 ;
        RECT 2.07 1.07 2.16 1.48 ;
        RECT 1.57 1.07 1.66 1.48 ;
        RECT 1.07 1.07 1.16 1.48 ;
        RECT 0.57 1.07 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.8 0.08 ;
        RECT 2.32 -0.08 2.41 0.345 ;
        RECT 1.795 -0.08 1.935 0.32 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.05 0.625 0.23 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.22 0.605 2.51 0.745 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.795 0.425 1.945 0.605 ;
      LAYER MET2 ;
        RECT 1.85 0.225 1.95 0.76 ;
      LAYER VIA1 ;
        RECT 1.855 0.455 1.945 0.545 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.79 0.89 1.935 0.98 ;
        RECT 1.055 0.33 1.145 0.98 ;
        RECT 0.795 0.33 1.145 0.42 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.04 0.84 2.435 0.93 ;
      RECT 2.04 0.33 2.13 0.93 ;
      RECT 1.255 0.695 2.13 0.785 ;
      RECT 1.255 0.635 1.545 0.785 ;
      RECT 2.04 0.33 2.185 0.42 ;
      RECT 0.32 0.305 0.41 0.95 ;
      RECT 0.32 0.66 0.865 0.75 ;
  END
END NAND3BBX4H7R

MACRO NAND3BBX6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BBX6H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.535 1.07 1.625 1.48 ;
        RECT 1.005 1.095 1.145 1.48 ;
        RECT 0.535 1.055 0.625 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.535 -0.08 1.625 0.33 ;
        RECT 0.51 -0.08 0.65 0.32 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.42 0.545 0.72 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.655 0.615 1.745 0.975 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.41 0.615 1.545 0.815 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.74 0.915 1.395 1.005 ;
        RECT 0.995 0.255 1.085 1.005 ;
        RECT 0.74 0.255 1.085 0.345 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.56 ;
      LAYER VIA1 ;
        RECT 0.855 0.255 0.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.76 1.065 1.925 1.155 ;
      RECT 1.835 0.435 1.925 1.155 ;
      RECT 1.18 0.435 1.27 0.705 ;
      RECT 1.18 0.435 1.925 0.525 ;
      RECT 1.785 0.33 1.875 0.525 ;
      RECT 0.26 0.85 0.584 0.94 ;
      RECT 0.26 0.85 0.63 0.917 ;
      RECT 0.546 0.831 0.676 0.871 ;
      RECT 0.26 0.255 0.35 0.94 ;
      RECT 0.584 0.789 0.676 0.871 ;
      RECT 0.63 0.743 0.722 0.825 ;
      RECT 0.676 0.697 0.768 0.779 ;
      RECT 0.676 0.697 0.799 0.741 ;
      RECT 0.811 0.585 0.905 0.725 ;
      RECT 0.722 0.651 0.905 0.725 ;
      RECT 0.799 0.591 0.905 0.725 ;
      RECT 0.768 0.612 0.905 0.725 ;
      RECT 0.26 0.255 0.4 0.345 ;
  END
END NAND3BBX6H7R

MACRO NAND3BX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BX0P5H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.81 1.185 0.95 1.48 ;
        RECT 0.32 1.05 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.4 0.605 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.595 0.425 0.82 0.545 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.655 1.02 0.795 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.11 0.23 1.2 1.135 ;
        RECT 0.545 1.005 1.2 1.095 ;
        RECT 1.025 0.23 1.2 0.345 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.56 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.205 0.16 1.135 ;
      RECT 0.07 0.745 0.56 0.835 ;
  END
END NAND3BX0P5H7R

MACRO NAND3BX0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BX0P7H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.84 1.155 0.98 1.48 ;
        RECT 0.335 1.05 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.335 -0.08 0.425 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.4 0.605 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.425 0.85 0.545 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.655 1.02 0.795 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.575 0.975 1.245 1.065 ;
        RECT 1.155 0.225 1.245 1.065 ;
        RECT 1.055 0.225 1.245 0.375 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.56 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.205 0.16 1.155 ;
      RECT 0.07 0.745 0.56 0.835 ;
  END
END NAND3BX0P7H7R

MACRO NAND3BX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BX1H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.86 1.07 0.95 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.32 -0.08 0.41 0.335 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.405 0.6 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.445 0.85 0.565 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.015 0.61 1.165 0.79 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.61 0.89 1.345 0.98 ;
        RECT 1.255 0.29 1.345 0.98 ;
        RECT 1.1 0.29 1.345 0.38 ;
        RECT 1.125 0.89 1.215 1.075 ;
        RECT 0.61 0.89 0.7 1.06 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.205 0.16 1.155 ;
      RECT 0.07 0.71 0.615 0.8 ;
  END
END NAND3BX1H7R

MACRO NAND3BX1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BX1P4H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.835 1.095 0.975 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.4 0.605 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.455 0.825 0.6 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.59 1.16 0.79 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.585 0.905 1.345 0.995 ;
        RECT 1.255 0.325 1.345 0.995 ;
        RECT 1.1 0.325 1.345 0.415 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.205 0.16 1.155 ;
      RECT 0.07 0.71 0.575 0.8 ;
  END
END NAND3BX1P4H7R

MACRO NAND3BX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BX2H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.835 1.07 0.925 1.48 ;
        RECT 0.335 1.07 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.36 0.825 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.55 0.775 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.945 0.625 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.6 1.15 1.135 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.585 0.865 1.325 0.955 ;
        RECT 1.235 0.255 1.325 0.955 ;
        RECT 0.99 0.255 1.325 0.345 ;
        RECT 1.085 0.865 1.175 1.18 ;
        RECT 0.585 0.865 0.675 1.21 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.385 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 1.04 0.2 1.13 ;
      RECT 0.045 0.205 0.135 1.13 ;
      RECT 0.455 0.445 0.545 0.705 ;
      RECT 0.045 0.445 0.545 0.535 ;
      RECT 0.045 0.205 0.16 0.535 ;
  END
END NAND3BX2H7R

MACRO NAND3BX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BX3H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 2.055 1.095 2.195 1.48 ;
        RECT 1.555 1.095 1.695 1.48 ;
        RECT 1.055 1.095 1.195 1.48 ;
        RECT 0.795 1.095 0.935 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 0.795 -0.08 0.935 0.305 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.805 0.405 0.955 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.205 0.655 1.545 0.745 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.705 0.655 2.045 0.745 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.545 0.915 2.345 1.005 ;
        RECT 2.255 0.425 2.345 1.005 ;
        RECT 1.805 0.425 2.345 0.515 ;
        RECT 1.805 0.915 1.945 1.02 ;
        RECT 1.805 0.35 1.945 0.515 ;
        RECT 1.305 0.915 1.445 1.02 ;
        RECT 0.545 0.915 0.685 1.02 ;
      LAYER MET2 ;
        RECT 2.25 0.63 2.35 1.16 ;
      LAYER VIA1 ;
        RECT 2.255 0.855 2.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.055 0.17 2.195 0.335 ;
      RECT 1.555 0.17 1.695 0.335 ;
      RECT 1.04 0.17 2.195 0.26 ;
      RECT 0.57 0.395 1.445 0.485 ;
      RECT 1.305 0.35 1.445 0.485 ;
      RECT 0.57 0.295 0.66 0.485 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 0.045 0.625 0.785 0.715 ;
      RECT 0.045 0.23 0.185 0.32 ;
  END
END NAND3BX3H7R

MACRO NAND3BX4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BX4H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 2.005 1.07 2.095 1.48 ;
        RECT 1.49 1.07 1.58 1.48 ;
        RECT 0.87 1.07 0.96 1.48 ;
        RECT 0.335 1.07 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 0.82 -0.08 0.91 0.345 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.63 0.405 0.78 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.145 0.655 1.485 0.745 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.655 0.625 1.96 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.595 0.885 2.145 0.975 ;
        RECT 2.055 0.395 2.145 0.975 ;
        RECT 1.775 0.395 2.145 0.485 ;
        RECT 1.74 0.885 1.83 1.2 ;
        RECT 1.24 0.885 1.33 1.2 ;
        RECT 0.595 0.885 0.71 1.2 ;
      LAYER MET2 ;
        RECT 2.05 0.63 2.15 1.16 ;
      LAYER VIA1 ;
        RECT 2.055 0.855 2.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.025 0.215 1.165 0.32 ;
      RECT 1.025 0.215 2.165 0.305 ;
      RECT 0.691 0.435 1.415 0.525 ;
      RECT 1.275 0.395 1.415 0.525 ;
      RECT 0.66 0.381 0.691 0.51 ;
      RECT 0.616 0.416 0.729 0.472 ;
      RECT 0.57 0.26 0.66 0.427 ;
      RECT 0.045 0.925 0.2 1.015 ;
      RECT 0.045 0.255 0.135 1.015 ;
      RECT 0.495 0.62 0.835 0.71 ;
      RECT 0.495 0.609 0.654 0.71 ;
      RECT 0.495 0.576 0.633 0.71 ;
      RECT 0.484 0.455 0.495 0.584 ;
      RECT 0.484 0.53 0.587 0.584 ;
      RECT 0.446 0.53 0.587 0.559 ;
      RECT 0.045 0.45 0.484 0.54 ;
      RECT 0.045 0.484 0.541 0.54 ;
      RECT 0.045 0.255 0.16 0.54 ;
  END
END NAND3BX4H7R

MACRO NAND3BX6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BX6H7R 0 0 ;
  SIZE 3.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.2 1.48 ;
        RECT 2.535 1.07 2.625 1.48 ;
        RECT 2.035 1.07 2.125 1.48 ;
        RECT 1.535 1.07 1.625 1.48 ;
        RECT 1.035 1.07 1.125 1.48 ;
        RECT 0.535 0.87 0.625 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.2 0.08 ;
        RECT 1.01 -0.08 1.15 0.305 ;
        RECT 0.535 -0.08 0.625 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.6 0.59 0.78 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.44 0.655 1.98 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.18 0.655 2.72 0.745 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.76 0.885 2.945 0.975 ;
        RECT 2.855 0.395 2.945 0.975 ;
        RECT 2.785 0.885 2.875 1.2 ;
        RECT 2.26 0.395 2.945 0.485 ;
        RECT 2.785 0.275 2.875 0.485 ;
        RECT 2.285 0.885 2.375 1.2 ;
        RECT 1.785 0.885 1.875 1.2 ;
        RECT 1.285 0.885 1.375 1.2 ;
        RECT 0.76 0.885 0.875 1.2 ;
      LAYER MET2 ;
        RECT 2.85 0.63 2.95 1.16 ;
      LAYER VIA1 ;
        RECT 2.855 0.855 2.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.866 0.395 1.9 0.485 ;
      RECT 0.831 0.395 1.9 0.468 ;
      RECT 0.785 0.26 0.875 0.427 ;
      RECT 0.785 0.38 0.904 0.427 ;
      RECT 0.26 0.845 0.375 1.185 ;
      RECT 0.26 0.305 0.35 1.185 ;
      RECT 0.69 0.62 1.23 0.71 ;
      RECT 0.69 0.599 0.869 0.71 ;
      RECT 0.69 0.556 0.828 0.71 ;
      RECT 0.669 0.43 0.69 0.559 ;
      RECT 0.669 0.51 0.782 0.559 ;
      RECT 0.631 0.51 0.782 0.529 ;
      RECT 0.26 0.42 0.669 0.51 ;
      RECT 0.26 0.464 0.736 0.51 ;
      RECT 0.26 0.305 0.375 0.51 ;
      RECT 1.51 0.215 2.65 0.305 ;
  END
END NAND3BX6H7R

MACRO NAND3X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X0P5H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.56 1.075 0.7 1.48 ;
        RECT 0.07 1.05 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.39 0.655 0.59 0.79 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.645 0.305 0.745 0.575 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.84 0.205 0.945 1.15 ;
        RECT 0.32 0.895 0.945 0.985 ;
        RECT 0.32 0.895 0.41 1.135 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
END NAND3X0P5H7R

MACRO NAND3X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X0P7H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.56 1.09 0.7 1.48 ;
        RECT 0.07 1.05 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.395 0.625 0.545 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.645 0.42 0.765 0.645 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.84 0.91 0.945 1.118 ;
        RECT 0.855 0.23 0.945 1.118 ;
        RECT 0.84 0.23 0.945 0.37 ;
        RECT 0.32 0.91 0.945 1 ;
        RECT 0.32 0.91 0.41 1.103 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
END NAND3X0P7H7R

MACRO NAND3X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X1H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.565 1.095 0.705 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.62 0.23 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.37 0.42 0.545 0.575 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.635 0.59 0.75 0.825 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.84 0.225 0.945 1.075 ;
        RECT 0.32 0.915 0.945 1.005 ;
        RECT 0.32 0.915 0.41 1.06 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
END NAND3X1H7R

MACRO NAND3X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X1P4H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.545 1.095 0.685 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.365 0.625 0.545 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.355 0.745 0.655 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.84 0.3 0.945 1.031 ;
        RECT 0.295 0.901 0.945 0.991 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
END NAND3X1P4H7R

MACRO NAND3X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X2H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.705 1.05 1.795 1.48 ;
        RECT 1.135 1.185 1.275 1.48 ;
        RECT 0.58 1.185 0.72 1.48 ;
        RECT 0.06 1.075 0.2 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 0.295 -0.08 0.435 0.41 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.775 0.535 0.865 ;
        RECT 0.055 0.775 0.145 0.975 ;
      LAYER MET2 ;
        RECT 0.05 0.625 0.15 1.16 ;
      LAYER VIA1 ;
        RECT 0.055 0.855 0.145 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.725 0.655 1.065 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.625 0.79 1.775 0.945 ;
        RECT 1.435 0.79 1.775 0.88 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.245 0.61 1.705 0.7 ;
        RECT 1.565 0.35 1.705 0.7 ;
        RECT 1.455 1.005 1.545 1.175 ;
        RECT 0.315 1.005 1.545 1.095 ;
        RECT 1.245 0.61 1.345 1.095 ;
      LAYER MET2 ;
        RECT 1.45 0.84 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.84 0.17 1.93 0.45 ;
      RECT 1.34 0.17 1.43 0.45 ;
      RECT 0.8 0.17 1.93 0.26 ;
      RECT 0.07 0.5 0.635 0.59 ;
      RECT 0.545 0.35 0.635 0.59 ;
      RECT 0.07 0.31 0.16 0.59 ;
      RECT 0.545 0.35 1.215 0.44 ;
  END
END NAND3X2H7R

MACRO NAND3X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X3H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.705 1.035 1.795 1.48 ;
        RECT 1.135 1.09 1.275 1.48 ;
        RECT 0.56 1.09 0.7 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 0.295 -0.08 0.435 0.335 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.195 0.655 0.535 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.725 0.655 1.065 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.445 0.655 1.785 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.315 0.425 1.93 0.515 ;
        RECT 1.84 0.31 1.93 0.515 ;
        RECT 0.295 0.91 1.57 1 ;
        RECT 1.315 0.35 1.455 0.515 ;
        RECT 1.315 0.35 1.454 0.524 ;
        RECT 1.315 0.35 1.437 0.555 ;
        RECT 1.255 0.563 1.345 1 ;
        RECT 1.301 0.533 1.391 0.601 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.565 0.17 1.705 0.335 ;
      RECT 0.8 0.17 0.94 0.335 ;
      RECT 0.8 0.17 1.705 0.26 ;
      RECT 0.07 0.425 1.195 0.515 ;
      RECT 1.055 0.35 1.195 0.515 ;
      RECT 0.57 0.325 0.66 0.515 ;
      RECT 0.07 0.31 0.16 0.515 ;
  END
END NAND3X3H7R

MACRO NAND3X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X4H7R 0 0 ;
  SIZE 3.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.6 1.48 ;
        RECT 3.39 1.095 3.53 1.48 ;
        RECT 2.89 1.095 3.03 1.48 ;
        RECT 2.2 1.095 2.34 1.48 ;
        RECT 1.635 1.095 1.775 1.48 ;
        RECT 1.105 1.095 1.245 1.48 ;
        RECT 0.575 1.095 0.715 1.48 ;
        RECT 0.045 1.08 0.185 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.6 0.08 ;
        RECT 0.84 -0.08 0.98 0.26 ;
        RECT 0.31 -0.08 0.45 0.26 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.275 0.655 1.015 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.335 0.655 2.075 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.225 0.72 3.35 0.81 ;
        RECT 2.225 0.655 2.375 0.81 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.325 0.915 3.545 1.005 ;
        RECT 3.455 0.31 3.545 1.005 ;
        RECT 2.465 0.5 3.545 0.59 ;
        RECT 3.44 0.31 3.545 0.59 ;
        RECT 3.14 0.915 3.28 1.155 ;
        RECT 2.915 0.35 3.055 0.59 ;
        RECT 2.64 0.915 2.78 1.155 ;
        RECT 2.465 0.35 2.555 0.59 ;
        RECT 2.415 0.35 2.555 0.44 ;
        RECT 1.905 0.915 2.045 1.155 ;
        RECT 1.385 0.915 1.525 1.155 ;
        RECT 0.825 0.915 0.965 1.155 ;
        RECT 0.325 0.915 0.465 1.155 ;
      LAYER MET2 ;
        RECT 3.45 0.625 3.55 1.16 ;
      LAYER VIA1 ;
        RECT 3.455 0.855 3.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 3.165 0.17 3.305 0.41 ;
      RECT 2.665 0.17 2.805 0.41 ;
      RECT 1.37 0.17 3.305 0.26 ;
      RECT 0.045 0.35 2.305 0.44 ;
      RECT 0.045 0.335 0.185 0.44 ;
  END
END NAND3X4H7R

MACRO NAND3X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X6H7R 0 0 ;
  SIZE 3 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3 1.48 ;
        RECT 2.285 1.07 2.375 1.48 ;
        RECT 1.785 1.07 1.875 1.48 ;
        RECT 1.285 1.07 1.375 1.48 ;
        RECT 0.785 1.07 0.875 1.48 ;
        RECT 0.285 1.055 0.375 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3 0.08 ;
        RECT 0.76 -0.08 0.9 0.305 ;
        RECT 0.285 -0.08 0.375 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.655 0.98 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.18 0.655 1.72 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.93 0.655 2.47 0.745 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.51 0.885 2.745 0.975 ;
        RECT 2.655 0.395 2.745 0.975 ;
        RECT 2.01 0.395 2.745 0.485 ;
      LAYER MET2 ;
        RECT 2.65 0.63 2.75 1.16 ;
      LAYER VIA1 ;
        RECT 2.655 0.855 2.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.255 0.215 2.4 0.305 ;
      RECT 0.51 0.395 1.65 0.485 ;
  END
END NAND3X6H7R

MACRO NAND3X8H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X8H7R 0 0 ;
  SIZE 4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4 1.48 ;
        RECT 3.52 1.08 3.66 1.48 ;
        RECT 3.045 1.07 3.135 1.48 ;
        RECT 2.285 1.07 2.375 1.48 ;
        RECT 1.785 1.07 1.875 1.48 ;
        RECT 1.285 1.07 1.375 1.48 ;
        RECT 0.785 1.07 0.875 1.48 ;
        RECT 0.285 1.055 0.375 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4 0.08 ;
        RECT 1.01 -0.08 1.15 0.305 ;
        RECT 0.51 -0.08 0.65 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.655 1.195 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.655 2.195 0.745 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.725 0.655 3.465 0.745 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.51 0.885 3.745 0.975 ;
        RECT 3.655 0.395 3.745 0.975 ;
        RECT 2.77 0.395 3.745 0.485 ;
      LAYER MET2 ;
        RECT 3.65 0.63 3.75 1.16 ;
      LAYER VIA1 ;
        RECT 3.655 0.855 3.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.285 0.395 2.4 0.485 ;
      RECT 0.285 0.315 0.375 0.485 ;
      RECT 1.51 0.215 3.66 0.305 ;
  END
END NAND3X8H7R

MACRO NAND4BBX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BBX0P5H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.815 1.055 1.905 1.48 ;
        RECT 1.295 1.095 1.435 1.48 ;
        RECT 0.795 1.095 0.935 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.82 -0.08 1.91 0.345 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.385 0.625 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.765 0.625 1.945 0.775 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.845 0.395 0.99 0.555 ;
        RECT 0.845 0.395 0.945 0.595 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.625 1.24 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.25 1.15 0.785 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.57 0.91 1.425 1 ;
        RECT 1.335 0.35 1.425 1 ;
        RECT 1.055 0.91 1.16 1.175 ;
        RECT 0.57 0.91 0.66 1.14 ;
      LAYER MET2 ;
        RECT 1.05 1.015 1.15 1.22 ;
      LAYER VIA1 ;
        RECT 1.055 1.055 1.145 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.565 0.17 1.655 1.155 ;
      RECT 0.66 0.17 0.75 0.555 ;
      RECT 0.66 0.17 1.655 0.26 ;
      RECT 0.07 0.205 0.16 1.16 ;
      RECT 0.07 0.73 0.585 0.82 ;
  END
END NAND4BBX0P5H7R

MACRO NAND4BBX0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BBX0P7H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.815 1.055 1.905 1.48 ;
        RECT 1.295 1.09 1.435 1.48 ;
        RECT 0.795 1.095 0.935 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.82 -0.08 1.91 0.345 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.385 0.625 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.745 0.625 1.945 0.775 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.425 1.035 0.555 ;
        RECT 0.855 0.425 0.945 0.595 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.655 1.245 0.795 ;
      LAYER MET2 ;
        RECT 1.05 0.25 1.15 0.785 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.57 0.91 1.425 1 ;
        RECT 1.335 0.35 1.425 1 ;
        RECT 1.285 0.35 1.425 0.44 ;
        RECT 1.055 0.91 1.16 1.175 ;
        RECT 0.57 0.91 0.66 1.108 ;
      LAYER MET2 ;
        RECT 1.05 1.015 1.15 1.22 ;
      LAYER VIA1 ;
        RECT 1.055 1.055 1.145 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.565 0.17 1.655 1.155 ;
      RECT 0.67 0.17 0.76 0.58 ;
      RECT 0.67 0.17 1.655 0.26 ;
      RECT 0.07 0.205 0.16 1.155 ;
      RECT 0.07 0.73 0.585 0.82 ;
  END
END NAND4BBX0P7H7R

MACRO NAND4BBX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BBX1H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.815 1.055 1.905 1.48 ;
        RECT 1.295 1.095 1.435 1.48 ;
        RECT 0.795 1.095 0.935 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.82 -0.08 1.91 0.345 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.415 0.385 0.615 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.765 0.625 1.945 0.775 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.425 1.045 0.565 ;
        RECT 0.855 0.425 0.945 0.575 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.655 1.245 0.815 ;
      LAYER MET2 ;
        RECT 1.05 0.25 1.15 0.785 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.345 0.35 1.435 1.005 ;
        RECT 0.616 0.917 1.435 1.005 ;
        RECT 0.621 0.915 1.435 1.005 ;
        RECT 1.295 0.35 1.435 0.44 ;
        RECT 1.055 0.915 1.16 1.175 ;
        RECT 0.57 0.943 0.66 1.17 ;
      LAYER MET2 ;
        RECT 1.05 1.015 1.15 1.22 ;
      LAYER VIA1 ;
        RECT 1.055 1.055 1.145 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.565 0.17 1.655 1.155 ;
      RECT 0.66 0.17 0.75 0.615 ;
      RECT 0.66 0.17 1.655 0.26 ;
      RECT 0.07 0.205 0.16 1.16 ;
      RECT 0.07 0.75 0.565 0.84 ;
  END
END NAND4BBX1H7R

MACRO NAND4BBX1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BBX1P4H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.835 1.055 1.925 1.48 ;
        RECT 1.305 1.08 1.445 1.48 ;
        RECT 0.82 1.07 0.91 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.84 -0.08 1.93 0.345 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.795 0.405 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.765 0.625 1.945 0.775 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.425 0.99 0.65 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.585 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.82 1.37 0.975 ;
        RECT 1.28 0.705 1.37 0.975 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.08 0.375 1.46 0.465 ;
        RECT 1.08 0.375 1.17 0.737 ;
        RECT 1.075 0.698 1.165 1.016 ;
        RECT 0.57 0.855 1.165 0.945 ;
        RECT 0.57 0.855 0.66 1.016 ;
      LAYER MET2 ;
        RECT 0.85 0.815 0.95 1.22 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.585 0.195 1.675 1.155 ;
      RECT 0.665 0.195 0.755 0.765 ;
      RECT 0.665 0.195 1.675 0.285 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 0.045 0.535 0.535 0.625 ;
      RECT 0.045 0.23 0.185 0.32 ;
  END
END NAND4BBX1P4H7R

MACRO NAND4BBX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BBX2H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.835 1.055 1.925 1.48 ;
        RECT 1.345 1.055 1.435 1.48 ;
        RECT 0.82 1.07 0.91 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.835 -0.08 1.925 0.345 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.77 0.375 0.95 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.765 0.625 1.945 0.775 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.64 1.035 0.775 ;
        RECT 0.855 0.61 0.945 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.165 0.455 1.255 0.705 ;
        RECT 1.025 0.455 1.255 0.545 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.545 0.865 1.435 0.955 ;
        RECT 1.345 0.355 1.435 0.955 ;
        RECT 1.225 0.855 1.435 0.955 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.585 0.175 1.675 1.155 ;
      RECT 0.67 0.175 0.76 0.75 ;
      RECT 0.67 0.175 1.675 0.265 ;
      RECT 0.045 1.045 0.185 1.135 ;
      RECT 0.045 0.23 0.135 1.135 ;
      RECT 0.045 0.59 0.55 0.68 ;
      RECT 0.045 0.23 0.185 0.32 ;
  END
END NAND4BBX2H7R

MACRO NAND4BBX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BBX3H7R 0 0 ;
  SIZE 3.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.6 1.48 ;
        RECT 3.14 1.055 3.23 1.48 ;
        RECT 2.625 1.07 2.715 1.48 ;
        RECT 2.02 1.225 2.16 1.48 ;
        RECT 1.44 1.225 1.58 1.48 ;
        RECT 0.825 1.095 0.965 1.48 ;
        RECT 0.35 1.07 0.44 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.6 0.08 ;
        RECT 1.43 -0.08 1.57 0.175 ;
        RECT 0.36 -0.08 0.45 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.425 0.39 0.625 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.425 0.655 1.725 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.5 0.655 2.84 0.745 ;
      LAYER MET2 ;
        RECT 2.65 0.43 2.75 0.96 ;
      LAYER VIA1 ;
        RECT 2.655 0.655 2.745 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.97 0.455 3.06 0.63 ;
        RECT 2.26 0.455 3.06 0.545 ;
        RECT 2.26 0.455 2.35 0.63 ;
      LAYER MET2 ;
        RECT 2.45 0.225 2.55 0.76 ;
      LAYER VIA1 ;
        RECT 2.455 0.455 2.545 0.545 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.045 0.855 3.255 0.945 ;
        RECT 3.165 0.29 3.255 0.945 ;
        RECT 3.115 0.29 3.255 0.38 ;
        RECT 2.89 0.855 2.98 1.045 ;
        RECT 2.36 0.855 2.45 1.045 ;
        RECT 1.12 1.045 2.135 1.135 ;
        RECT 2.045 0.35 2.135 1.135 ;
        RECT 1.044 1.041 1.174 1.066 ;
        RECT 1.044 1.014 1.166 1.066 ;
        RECT 1.006 0.976 1.12 1.024 ;
        RECT 1.09 1.045 2.135 1.104 ;
        RECT 0.57 0.938 1.09 1.005 ;
        RECT 0.57 0.915 1.044 1.005 ;
        RECT 0.57 0.915 0.72 1.02 ;
      LAYER MET2 ;
        RECT 3.05 0.63 3.15 1.16 ;
      LAYER VIA1 ;
        RECT 3.055 0.855 3.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.855 0.265 1.684 0.355 ;
      RECT 2.625 0.17 2.715 0.33 ;
      RECT 0.855 0.265 1.752 0.31 ;
      RECT 1.611 0.242 1.779 0.274 ;
      RECT 1.684 0.181 1.706 0.344 ;
      RECT 1.706 0.17 2.715 0.26 ;
      RECT 1.657 0.205 2.715 0.26 ;
      RECT 1.291 0.865 1.93 0.955 ;
      RECT 1.84 0.355 1.93 0.955 ;
      RECT 1.288 0.825 1.291 0.954 ;
      RECT 1.242 0.801 1.288 0.929 ;
      RECT 1.196 0.755 1.242 0.883 ;
      RECT 1.196 0.846 1.329 0.883 ;
      RECT 1.15 0.709 1.196 0.837 ;
      RECT 1.104 0.663 1.15 0.791 ;
      RECT 1.066 0.709 1.196 0.749 ;
      RECT 0.75 0.64 1.104 0.73 ;
      RECT 1.815 0.355 1.93 0.495 ;
      RECT 0.07 1.04 0.215 1.13 ;
      RECT 0.07 0.23 0.16 1.13 ;
      RECT 0.07 0.715 0.59 0.805 ;
      RECT 0.5 0.455 0.59 0.805 ;
      RECT 0.07 0.23 0.165 0.805 ;
      RECT 1.24 0.455 1.33 0.63 ;
      RECT 0.5 0.455 1.33 0.545 ;
      RECT 0.07 0.23 0.21 0.32 ;
  END
END NAND4BBX3H7R

MACRO NAND4BBX4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BBX4H7R 0 0 ;
  SIZE 3.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.6 1.48 ;
        RECT 3.14 1.055 3.23 1.48 ;
        RECT 2.625 1.07 2.715 1.48 ;
        RECT 2.02 1.21 2.16 1.48 ;
        RECT 1.44 1.21 1.58 1.48 ;
        RECT 0.85 1.07 0.94 1.48 ;
        RECT 0.35 1.07 0.44 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.6 0.08 ;
        RECT 1.43 -0.08 1.57 0.175 ;
        RECT 0.36 -0.08 0.45 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.425 0.355 0.695 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.425 0.655 1.725 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.485 0.655 2.825 0.745 ;
      LAYER MET2 ;
        RECT 2.65 0.43 2.75 0.96 ;
      LAYER VIA1 ;
        RECT 2.655 0.655 2.745 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.985 0.539 3.075 0.705 ;
        RECT 2.25 0.494 3.031 0.545 ;
        RECT 2.25 0.463 2.985 0.545 ;
        RECT 2.969 0.539 3.075 0.591 ;
        RECT 2.25 0.455 2.969 0.545 ;
        RECT 2.931 0.539 3.075 0.564 ;
        RECT 2.25 0.455 2.34 0.705 ;
      LAYER MET2 ;
        RECT 2.45 0.225 2.55 0.76 ;
      LAYER VIA1 ;
        RECT 2.455 0.455 2.545 0.545 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.045 0.855 3.255 0.945 ;
        RECT 3.165 0.38 3.255 0.945 ;
        RECT 3.115 0.38 3.255 0.47 ;
        RECT 1.121 1.03 2.135 1.12 ;
        RECT 2.045 0.355 2.135 1.12 ;
        RECT 1.019 1.011 1.159 1.041 ;
        RECT 1.019 0.987 1.121 1.041 ;
        RECT 1.111 1.03 2.135 1.115 ;
        RECT 0.981 0.959 1.111 0.999 ;
        RECT 1.065 1.03 2.135 1.087 ;
        RECT 0.575 0.913 1.065 0.98 ;
        RECT 0.575 0.89 1.019 0.98 ;
      LAYER MET2 ;
        RECT 3.05 0.63 3.15 1.16 ;
      LAYER VIA1 ;
        RECT 3.055 0.855 3.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.87 0.265 1.684 0.355 ;
      RECT 2.625 0.17 2.715 0.33 ;
      RECT 0.87 0.265 1.752 0.31 ;
      RECT 1.611 0.242 1.779 0.274 ;
      RECT 1.684 0.181 1.706 0.344 ;
      RECT 1.706 0.17 2.715 0.26 ;
      RECT 1.657 0.205 2.715 0.26 ;
      RECT 1.222 0.85 1.91 0.94 ;
      RECT 1.82 0.355 1.91 0.94 ;
      RECT 1.213 0.807 1.222 0.936 ;
      RECT 1.167 0.78 1.213 0.908 ;
      RECT 1.121 0.734 1.167 0.862 ;
      RECT 1.121 0.831 1.26 0.862 ;
      RECT 1.075 0.688 1.121 0.816 ;
      RECT 1.037 0.734 1.167 0.774 ;
      RECT 0.735 0.665 1.075 0.755 ;
      RECT 1.815 0.355 1.91 0.495 ;
      RECT 0.07 0.815 0.215 1.01 ;
      RECT 0.07 0.815 0.404 0.905 ;
      RECT 0.07 0.815 0.45 0.882 ;
      RECT 0.366 0.796 0.496 0.836 ;
      RECT 0.07 0.23 0.165 1.01 ;
      RECT 0.404 0.754 0.5 0.811 ;
      RECT 0.45 0.708 0.546 0.786 ;
      RECT 0.496 0.683 0.5 0.811 ;
      RECT 0.5 0.455 0.59 0.741 ;
      RECT 1.245 0.455 1.335 0.705 ;
      RECT 0.5 0.455 1.335 0.545 ;
      RECT 0.07 0.23 0.21 0.32 ;
  END
END NAND4BBX4H7R

MACRO NAND4BBX6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BBX6H7R 0 0 ;
  SIZE 4.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.8 1.48 ;
        RECT 4.34 1.07 4.43 1.48 ;
        RECT 3.84 1.07 3.93 1.48 ;
        RECT 3.34 1.07 3.43 1.48 ;
        RECT 2.84 1.07 2.93 1.48 ;
        RECT 2.34 1.07 2.43 1.48 ;
        RECT 1.71 1.07 1.8 1.48 ;
        RECT 1.12 1.21 1.26 1.48 ;
        RECT 0.535 1.07 0.625 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.8 0.08 ;
        RECT 1.75 -0.08 1.89 0.2 ;
        RECT 1.18 -0.08 1.27 0.345 ;
        RECT 0.535 -0.08 0.625 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.425 0.545 0.725 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.645 0.595 0.795 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.995 0.655 3.535 0.745 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.735 0.655 4.275 0.745 ;
      LAYER MET2 ;
        RECT 3.85 0.43 3.95 0.96 ;
      LAYER VIA1 ;
        RECT 3.855 0.655 3.945 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.435 0.885 4.545 0.975 ;
        RECT 4.455 0.215 4.545 0.975 ;
        RECT 3.815 0.215 4.545 0.305 ;
      LAYER MET2 ;
        RECT 4.45 0.625 4.55 1.16 ;
      LAYER VIA1 ;
        RECT 4.455 0.855 4.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.885 0.85 1.025 0.94 ;
      RECT 0.885 0.355 0.975 0.94 ;
      RECT 1.87 0.625 2.785 0.715 ;
      RECT 1.87 0.47 1.96 0.715 ;
      RECT 0.885 0.47 1.96 0.56 ;
      RECT 2.09 0.395 2.705 0.485 ;
      RECT 2.09 0.29 2.18 0.485 ;
      RECT 1.435 0.29 2.18 0.38 ;
      RECT 0.806 1.03 1.22 1.12 ;
      RECT 1.13 0.655 1.22 1.12 ;
      RECT 0.771 0.974 0.806 1.103 ;
      RECT 0.725 0.934 0.771 1.062 ;
      RECT 0.725 1.011 0.844 1.062 ;
      RECT 0.679 0.888 0.725 1.016 ;
      RECT 0.641 0.865 0.679 0.974 ;
      RECT 0.26 0.865 0.679 0.955 ;
      RECT 0.26 0.24 0.35 0.955 ;
      RECT 1.13 0.655 1.71 0.745 ;
      RECT 0.26 0.24 0.375 0.38 ;
      RECT 3.065 0.395 4.205 0.485 ;
      RECT 2.315 0.215 3.455 0.305 ;
  END
END NAND4BBX6H7R

MACRO NAND4BX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BX0P5H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.37 1.1 1.51 1.48 ;
        RECT 0.84 1.1 0.98 1.48 ;
        RECT 0.335 1.05 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.335 -0.08 0.425 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.4 0.605 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.61 0.455 0.88 0.555 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.655 1.125 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.545 1.355 0.815 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.6 0.92 1.545 1.01 ;
        RECT 1.455 0.23 1.545 1.01 ;
        RECT 1.355 0.23 1.545 0.32 ;
        RECT 1.13 0.92 1.22 1.12 ;
        RECT 0.6 0.92 0.69 1.12 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.205 0.16 1.13 ;
      RECT 0.07 0.74 0.56 0.83 ;
  END
END NAND4BX0P5H7R

MACRO NAND4BX0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BX0P7H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.325 1.06 1.465 1.48 ;
        RECT 0.825 1.075 0.965 1.48 ;
        RECT 0.335 1.05 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.335 -0.08 0.425 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.4 0.605 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.58 0.455 0.88 0.545 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.655 1.095 0.755 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.52 1.355 0.79 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.6 0.88 1.545 0.97 ;
        RECT 1.455 0.255 1.545 0.97 ;
        RECT 1.325 0.255 1.545 0.345 ;
        RECT 1.1 0.88 1.19 1.09 ;
        RECT 0.6 0.88 0.69 1.09 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.205 0.16 1.135 ;
      RECT 0.07 0.705 0.56 0.795 ;
  END
END NAND4BX0P7H7R

MACRO NAND4BX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BX1H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.37 1.11 1.51 1.48 ;
        RECT 0.84 1.11 0.98 1.48 ;
        RECT 0.335 1.04 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.335 -0.08 0.425 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.4 0.605 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.625 0.8 0.815 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.425 1.145 0.575 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.245 0.61 1.365 0.835 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.575 0.93 1.545 1.02 ;
        RECT 1.455 0.28 1.545 1.02 ;
        RECT 1.355 0.28 1.545 0.37 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.205 0.16 1.125 ;
      RECT 0.07 0.735 0.565 0.825 ;
  END
END NAND4BX1H7R

MACRO NAND4BX1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BX1P4H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.355 1.065 1.495 1.48 ;
        RECT 0.84 1.065 0.98 1.48 ;
        RECT 0.335 1.04 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.335 -0.08 0.425 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.4 0.605 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.75 0.455 0.84 0.65 ;
        RECT 0.625 0.455 0.84 0.545 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.425 1.145 0.65 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.245 0.55 1.365 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.6 0.885 1.545 0.975 ;
        RECT 1.455 0.325 1.545 0.975 ;
        RECT 1.355 0.325 1.545 0.415 ;
        RECT 0.6 0.885 0.69 1.025 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.205 0.16 1.125 ;
      RECT 0.07 0.7 0.605 0.79 ;
  END
END NAND4BX1P4H7R

MACRO NAND4BX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BX2H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.495 1.055 1.585 1.48 ;
        RECT 0.995 1.07 1.085 1.48 ;
        RECT 0.485 0.87 0.575 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 0.535 -0.08 0.625 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.365 0.625 0.545 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.425 0.955 0.705 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.595 1.205 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.365 0.625 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.605 1.55 1.135 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.72 0.87 1.725 0.96 ;
        RECT 1.635 0.255 1.725 0.96 ;
        RECT 1.4 0.255 1.725 0.345 ;
      LAYER MET2 ;
        RECT 1.45 0.18 1.55 0.385 ;
      LAYER VIA1 ;
        RECT 1.455 0.255 1.545 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.185 0.865 0.35 1.155 ;
      RECT 0.185 0.445 0.275 1.155 ;
      RECT 0.635 0.445 0.725 0.705 ;
      RECT 0.185 0.445 0.725 0.535 ;
      RECT 0.285 0.31 0.375 0.535 ;
  END
END NAND4BX2H7R

MACRO NAND4BX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BX3H7R 0 0 ;
  SIZE 3 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3 1.48 ;
        RECT 2.755 1.095 2.895 1.48 ;
        RECT 2.055 1.095 2.195 1.48 ;
        RECT 1.555 1.095 1.695 1.48 ;
        RECT 1.055 1.095 1.195 1.48 ;
        RECT 0.795 1.095 0.935 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3 0.08 ;
        RECT 0.795 -0.08 0.935 0.305 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.8 0.405 0.95 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.205 0.655 1.545 0.745 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.705 0.655 2.045 0.745 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.46 0.625 2.75 0.775 ;
      LAYER MET2 ;
        RECT 2.65 0.43 2.75 0.96 ;
      LAYER VIA1 ;
        RECT 2.655 0.655 2.745 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.545 0.915 2.945 1.005 ;
        RECT 2.84 0.17 2.945 1.005 ;
        RECT 2.315 0.17 2.945 0.26 ;
        RECT 2.505 0.915 2.645 1.02 ;
        RECT 2.315 0.17 2.455 0.335 ;
        RECT 1.805 0.915 1.945 1.02 ;
        RECT 1.305 0.915 1.445 1.02 ;
        RECT 0.545 0.915 0.685 1.02 ;
      LAYER MET2 ;
        RECT 2.85 0.63 2.95 1.16 ;
      LAYER VIA1 ;
        RECT 2.855 0.855 2.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.805 0.425 2.705 0.515 ;
      RECT 2.565 0.35 2.705 0.515 ;
      RECT 1.805 0.35 1.945 0.515 ;
      RECT 1.58 0.17 1.67 0.36 ;
      RECT 2.055 0.17 2.195 0.335 ;
      RECT 1.04 0.17 2.195 0.26 ;
      RECT 0.545 0.395 1.445 0.485 ;
      RECT 1.305 0.35 1.445 0.485 ;
      RECT 0.545 0.315 0.685 0.485 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 0.045 0.61 0.785 0.7 ;
      RECT 0.045 0.23 0.185 0.32 ;
  END
END NAND4BX3H7R

MACRO NAND4BX4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BX4H7R 0 0 ;
  SIZE 3.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.2 1.48 ;
        RECT 2.72 1.07 2.81 1.48 ;
        RECT 2.005 1.07 2.095 1.48 ;
        RECT 1.49 1.07 1.58 1.48 ;
        RECT 0.87 1.07 0.96 1.48 ;
        RECT 0.335 1.07 0.425 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.2 0.08 ;
        RECT 0.795 -0.08 0.935 0.32 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.24 0.605 0.36 0.83 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.145 0.655 1.485 0.745 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.645 0.655 1.985 0.745 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.375 0.655 2.715 0.745 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.595 0.885 2.945 0.975 ;
        RECT 2.855 0.215 2.945 0.975 ;
        RECT 2.76 0.215 2.945 0.32 ;
        RECT 2.255 0.215 2.945 0.305 ;
        RECT 2.47 0.885 2.56 1.2 ;
        RECT 2.255 0.215 2.395 0.32 ;
        RECT 1.74 0.885 1.83 1.2 ;
        RECT 1.24 0.885 1.33 1.2 ;
        RECT 0.595 0.885 0.685 1.2 ;
      LAYER MET2 ;
        RECT 2.85 0.63 2.95 1.16 ;
      LAYER VIA1 ;
        RECT 2.855 0.855 2.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.775 0.41 2.645 0.5 ;
      RECT 2.505 0.395 2.645 0.5 ;
      RECT 1.775 0.395 1.915 0.5 ;
      RECT 2.025 0.215 2.165 0.32 ;
      RECT 1.025 0.215 1.165 0.32 ;
      RECT 1.025 0.215 2.165 0.305 ;
      RECT 0.646 0.41 1.415 0.5 ;
      RECT 1.275 0.395 1.415 0.5 ;
      RECT 0.616 0.41 1.415 0.485 ;
      RECT 0.57 0.284 0.66 0.447 ;
      RECT 0.57 0.398 0.684 0.447 ;
      RECT 0.06 0.92 0.2 1.01 ;
      RECT 0.06 0.305 0.15 1.01 ;
      RECT 0.495 0.62 0.835 0.71 ;
      RECT 0.495 0.619 0.634 0.71 ;
      RECT 0.495 0.596 0.633 0.71 ;
      RECT 0.485 0.476 0.495 0.604 ;
      RECT 0.485 0.55 0.587 0.604 ;
      RECT 0.439 0.448 0.485 0.576 ;
      RECT 0.439 0.504 0.541 0.576 ;
      RECT 0.401 0.504 0.541 0.534 ;
      RECT 0.06 0.425 0.439 0.515 ;
      RECT 0.06 0.305 0.16 0.515 ;
  END
END NAND4BX4H7R

MACRO NAND4BX6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BX6H7R 0 0 ;
  SIZE 4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4 1.48 ;
        RECT 3.51 1.08 3.65 1.48 ;
        RECT 3.035 1.07 3.125 1.48 ;
        RECT 2.535 1.07 2.625 1.48 ;
        RECT 2.035 1.07 2.125 1.48 ;
        RECT 1.535 1.07 1.625 1.48 ;
        RECT 1.035 1.07 1.125 1.48 ;
        RECT 0.535 0.87 0.625 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4 0.08 ;
        RECT 1.01 -0.08 1.15 0.305 ;
        RECT 0.535 -0.08 0.625 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.6 0.59 0.78 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.44 0.655 1.98 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.18 0.655 2.72 0.745 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.905 0.655 3.445 0.745 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.76 0.885 3.625 0.975 ;
        RECT 3.535 0.215 3.625 0.975 ;
        RECT 3.425 0.855 3.625 0.975 ;
        RECT 3.01 0.215 3.625 0.305 ;
        RECT 3.285 0.885 3.375 1.2 ;
        RECT 2.785 0.885 2.875 1.2 ;
        RECT 2.285 0.885 2.375 1.2 ;
        RECT 1.785 0.885 1.875 1.2 ;
        RECT 1.285 0.885 1.375 1.2 ;
        RECT 0.76 0.885 0.9 1.175 ;
      LAYER MET2 ;
        RECT 3.45 0.625 3.55 1.16 ;
      LAYER VIA1 ;
        RECT 3.455 0.855 3.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.866 0.395 1.9 0.485 ;
      RECT 0.831 0.395 1.9 0.468 ;
      RECT 0.785 0.26 0.875 0.427 ;
      RECT 0.785 0.38 0.904 0.427 ;
      RECT 0.26 0.88 0.4 1.17 ;
      RECT 0.26 0.305 0.35 1.17 ;
      RECT 0.69 0.62 1.23 0.71 ;
      RECT 0.69 0.599 0.869 0.71 ;
      RECT 0.69 0.556 0.828 0.71 ;
      RECT 0.669 0.43 0.69 0.559 ;
      RECT 0.669 0.51 0.782 0.559 ;
      RECT 0.631 0.51 0.782 0.529 ;
      RECT 0.26 0.42 0.669 0.51 ;
      RECT 0.26 0.464 0.736 0.51 ;
      RECT 0.26 0.305 0.375 0.51 ;
      RECT 2.26 0.395 3.4 0.485 ;
      RECT 1.51 0.215 2.65 0.305 ;
  END
END NAND4BX6H7R

MACRO NAND4X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X0P5H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.855 1.03 0.995 1.48 ;
        RECT 0.325 1.03 0.465 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.085 -0.08 0.175 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.15 0.635 0.375 0.755 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.385 0.425 0.61 0.545 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.635 0.85 0.755 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.425 1.145 0.65 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.085 0.85 1.345 0.94 ;
        RECT 1.255 0.23 1.345 0.94 ;
        RECT 1.12 0.23 1.345 0.32 ;
        RECT 1.145 0.85 1.235 1.09 ;
        RECT 0.615 0.85 0.705 1.075 ;
        RECT 0.085 0.85 0.175 1.09 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END Y
END NAND4X0P5H7R

MACRO NAND4X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X0P7H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.855 1.03 0.995 1.48 ;
        RECT 0.325 1.03 0.465 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.085 -0.08 0.175 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.15 0.64 0.375 0.76 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.385 0.425 0.61 0.545 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.64 0.85 0.76 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.425 1.145 0.65 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.085 0.85 1.345 0.94 ;
        RECT 1.255 0.245 1.345 0.94 ;
        RECT 1.12 0.245 1.345 0.335 ;
        RECT 1.145 0.85 1.235 1.058 ;
        RECT 0.615 0.85 0.705 1.043 ;
        RECT 0.085 0.85 0.175 1.058 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END Y
END NAND4X0P7H7R

MACRO NAND4X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X1H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.855 1.05 0.995 1.48 ;
        RECT 0.325 1.05 0.465 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.085 -0.08 0.175 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.075 0.655 0.375 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.37 0.445 0.595 0.565 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.655 0.85 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.625 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.06 0.87 1.345 0.96 ;
        RECT 1.255 0.29 1.345 0.96 ;
        RECT 1.12 0.29 1.345 0.38 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END Y
END NAND4X1H7R

MACRO NAND4X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X1P4H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.855 1.05 0.995 1.48 ;
        RECT 0.325 1.05 0.465 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.085 -0.08 0.175 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.435 0.425 0.555 0.65 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.595 0.805 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.425 1.145 0.65 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.085 0.87 1.345 0.96 ;
        RECT 1.255 0.245 1.345 0.96 ;
        RECT 1.12 0.245 1.345 0.335 ;
        RECT 0.085 0.87 0.175 1.01 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END Y
END NAND4X1P4H7R

MACRO NAND4X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X2H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.995 1.07 1.085 1.48 ;
        RECT 0.495 1.07 0.585 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.285 -0.08 0.375 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.2 0.645 0.47 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.595 0.595 0.745 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.405 0.945 0.705 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.045 0.595 1.195 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.22 0.865 1.375 0.955 ;
        RECT 1.285 0.255 1.375 0.955 ;
        RECT 1.185 0.255 1.375 0.345 ;
      LAYER MET2 ;
        RECT 1.25 0.18 1.35 0.56 ;
      LAYER VIA1 ;
        RECT 1.255 0.255 1.345 0.345 ;
    END
  END Y
END NAND4X2H7R

MACRO NAND4X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X3H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 2.3 1.055 2.39 1.48 ;
        RECT 1.77 1.07 1.86 1.48 ;
        RECT 1.14 1.07 1.23 1.48 ;
        RECT 0.57 1.07 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.195 0.655 0.535 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.725 0.655 1.065 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.425 0.655 1.765 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.925 0.655 2.265 0.745 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.32 0.855 2.445 0.945 ;
        RECT 2.355 0.395 2.445 0.945 ;
        RECT 2.07 0.395 2.445 0.485 ;
        RECT 2.07 0.35 2.21 0.485 ;
        RECT 2.05 0.855 2.14 1.045 ;
        RECT 1.52 0.855 1.61 1.045 ;
        RECT 0.85 0.855 0.94 1.045 ;
        RECT 0.32 0.855 0.41 1.045 ;
      LAYER MET2 ;
        RECT 2.25 0.63 2.35 1.16 ;
      LAYER VIA1 ;
        RECT 2.255 0.855 2.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.29 0.395 1.92 0.485 ;
      RECT 1.83 0.17 1.92 0.485 ;
      RECT 1.29 0.35 1.43 0.485 ;
      RECT 2.335 0.17 2.475 0.305 ;
      RECT 1.83 0.17 2.475 0.26 ;
      RECT 1.555 0.17 1.695 0.305 ;
      RECT 0.795 0.17 0.935 0.305 ;
      RECT 0.795 0.17 1.695 0.26 ;
      RECT 0.07 0.395 1.2 0.485 ;
      RECT 1.06 0.35 1.2 0.485 ;
      RECT 0.57 0.295 0.66 0.485 ;
      RECT 0.07 0.28 0.16 0.485 ;
  END
END NAND4X3H7R

MACRO NAND4X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X4H7R 0 0 ;
  SIZE 3 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3 1.48 ;
        RECT 2.52 1.07 2.61 1.48 ;
        RECT 1.96 1.07 2.05 1.48 ;
        RECT 1.36 1.07 1.45 1.48 ;
        RECT 0.79 1.07 0.88 1.48 ;
        RECT 0.29 1.055 0.38 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3 0.08 ;
        RECT 0.515 -0.08 0.655 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.415 0.635 0.755 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.945 0.655 1.285 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.615 0.655 1.955 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.115 0.655 2.455 0.745 ;
      LAYER MET2 ;
        RECT 2.25 0.255 2.35 0.785 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.515 0.885 2.815 0.975 ;
        RECT 2.725 0.215 2.815 0.975 ;
        RECT 2.245 0.215 2.815 0.305 ;
        RECT 2.255 0.885 2.345 1.2 ;
        RECT 1.71 0.885 1.8 1.2 ;
        RECT 1.07 0.885 1.16 1.2 ;
        RECT 0.515 0.885 0.63 1.2 ;
      LAYER MET2 ;
        RECT 2.25 1.015 2.35 1.22 ;
      LAYER VIA1 ;
        RECT 2.255 1.055 2.345 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.495 0.395 2.635 0.485 ;
      RECT 1.495 0.38 1.635 0.485 ;
      RECT 1.745 0.19 1.885 0.305 ;
      RECT 1.015 0.19 1.155 0.305 ;
      RECT 1.015 0.19 1.885 0.28 ;
      RECT 0.29 0.395 1.405 0.485 ;
      RECT 1.265 0.38 1.405 0.485 ;
      RECT 0.29 0.305 0.38 0.485 ;
  END
END NAND4X4H7R

MACRO NAND4X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X6H7R 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.8 1.48 ;
        RECT 3.325 1.07 3.415 1.48 ;
        RECT 2.825 1.07 2.915 1.48 ;
        RECT 2.325 1.07 2.415 1.48 ;
        RECT 1.825 1.07 1.915 1.48 ;
        RECT 1.325 1.07 1.415 1.48 ;
        RECT 0.825 1.07 0.915 1.48 ;
        RECT 0.325 1.055 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.8 0.08 ;
        RECT 0.8 -0.08 0.94 0.305 ;
        RECT 0.325 -0.08 0.415 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.48 0.655 1.02 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.22 0.655 1.76 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.97 0.655 2.51 0.745 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.72 0.655 3.26 0.745 ;
      LAYER MET2 ;
        RECT 2.85 0.43 2.95 0.96 ;
      LAYER VIA1 ;
        RECT 2.855 0.655 2.945 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 0.885 3.545 0.975 ;
        RECT 3.455 0.215 3.545 0.975 ;
        RECT 2.8 0.215 3.545 0.305 ;
      LAYER MET2 ;
        RECT 3.45 0.625 3.55 1.16 ;
      LAYER VIA1 ;
        RECT 3.455 0.855 3.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.05 0.395 3.19 0.485 ;
      RECT 1.3 0.215 2.44 0.305 ;
      RECT 0.55 0.395 1.69 0.485 ;
  END
END NAND4X6H7R

MACRO NOR2BX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BX0P5H7R 0 0 ;
  SIZE 1.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.2 1.48 ;
        RECT 0.375 0.895 0.465 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.2 0.08 ;
        RECT 0.92 -0.08 1.06 0.175 ;
        RECT 0.375 -0.08 0.465 0.35 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.625 0.4 0.805 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.625 0.835 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.945 0.825 1.145 0.98 ;
        RECT 0.945 0.265 1.035 0.98 ;
        RECT 0.65 0.265 1.035 0.355 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END Z
  OBS
    LAYER MET1 ;
      RECT 0.07 0.225 0.16 0.98 ;
      RECT 0.07 0.445 0.615 0.535 ;
  END
END NOR2BX0P5H7R

MACRO NOR2BX0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BX0P7H7R 0 0 ;
  SIZE 1.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.2 1.48 ;
        RECT 0.375 0.895 0.465 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.2 0.08 ;
        RECT 0.92 -0.08 1.06 0.175 ;
        RECT 0.375 -0.08 0.465 0.35 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.625 0.4 0.805 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.64 0.835 0.78 ;
      LAYER MET2 ;
        RECT 0.65 0.6 0.75 1.135 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.925 0.265 1.015 0.98 ;
        RECT 0.625 0.265 1.015 0.355 ;
        RECT 0.625 0.255 0.775 0.355 ;
      LAYER MET2 ;
        RECT 0.65 0.18 0.75 0.385 ;
      LAYER VIA1 ;
        RECT 0.655 0.255 0.745 0.345 ;
    END
  END Z
  OBS
    LAYER MET1 ;
      RECT 0.07 0.215 0.16 0.98 ;
      RECT 0.475 0.445 0.615 0.55 ;
      RECT 0.07 0.445 0.615 0.535 ;
  END
END NOR2BX0P7H7R

MACRO NOR2BX12H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BX12H7R 0 0 ;
  SIZE 4.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.2 1.48 ;
        RECT 2.21 1.08 2.35 1.48 ;
        RECT 1.71 1.095 1.85 1.48 ;
        RECT 1.21 1.095 1.35 1.48 ;
        RECT 0.72 1.07 0.81 1.48 ;
        RECT 0.22 1.055 0.31 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.2 0.08 ;
        RECT 3.757 -0.08 3.897 0.305 ;
        RECT 3.257 -0.08 3.397 0.305 ;
        RECT 2.757 -0.08 2.897 0.305 ;
        RECT 2.257 -0.08 2.397 0.305 ;
        RECT 1.757 -0.08 1.897 0.305 ;
        RECT 1.257 -0.08 1.397 0.305 ;
        RECT 0.757 -0.08 0.897 0.305 ;
        RECT 0.282 -0.08 0.372 0.345 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.65 0.615 0.77 0.84 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.625 0.655 3.765 0.745 ;
      LAYER MET2 ;
        RECT 2.85 0.43 2.95 0.96 ;
      LAYER VIA1 ;
        RECT 2.855 0.655 2.945 0.745 ;
    END
  END B
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.69 0.885 3.945 0.975 ;
        RECT 3.855 0.395 3.945 0.975 ;
        RECT 1.057 0.395 3.945 0.485 ;
        RECT 1.057 0.235 1.147 0.485 ;
        RECT 1.007 0.235 1.147 0.325 ;
      LAYER MET2 ;
        RECT 3.85 0.43 3.95 0.96 ;
      LAYER VIA1 ;
        RECT 3.855 0.655 3.945 0.745 ;
    END
  END Z
  OBS
    LAYER MET1 ;
      RECT 2.49 1.065 4.08 1.155 ;
      RECT 2.49 0.9 2.58 1.155 ;
      RECT 0.96 0.9 2.58 0.99 ;
      RECT 0.47 0.395 0.56 0.95 ;
      RECT 0.86 0.64 2.03 0.73 ;
      RECT 0.86 0.395 0.95 0.73 ;
      RECT 0.47 0.395 0.95 0.485 ;
  END
END NOR2BX12H7R

MACRO NOR2BX16H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BX16H7R 0 0 ;
  SIZE 5.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.6 1.48 ;
        RECT 3.01 1.08 3.15 1.48 ;
        RECT 2.51 1.095 2.65 1.48 ;
        RECT 2.01 1.095 2.15 1.48 ;
        RECT 1.51 1.095 1.65 1.48 ;
        RECT 1.035 1.07 1.125 1.48 ;
        RECT 0.535 1.07 0.625 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.6 0.08 ;
        RECT 5.01 -0.08 5.15 0.305 ;
        RECT 4.51 -0.08 4.65 0.305 ;
        RECT 4.01 -0.08 4.15 0.305 ;
        RECT 3.51 -0.08 3.65 0.305 ;
        RECT 3.01 -0.08 3.15 0.305 ;
        RECT 2.51 -0.08 2.65 0.305 ;
        RECT 2.01 -0.08 2.15 0.305 ;
        RECT 1.51 -0.08 1.65 0.305 ;
        RECT 1.01 -0.08 1.15 0.305 ;
        RECT 0.51 -0.08 0.65 0.305 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.935 0.825 1.145 0.975 ;
        RECT 0.935 0.615 1.025 0.975 ;
        RECT 0.51 0.64 1.025 0.73 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.19 0.655 4.93 0.745 ;
      LAYER MET2 ;
        RECT 3.65 0.43 3.75 0.96 ;
      LAYER VIA1 ;
        RECT 3.655 0.655 3.745 0.745 ;
    END
  END B
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.49 0.885 5.145 0.975 ;
        RECT 5.055 0.395 5.145 0.975 ;
        RECT 1.31 0.395 5.145 0.485 ;
        RECT 1.31 0.215 1.4 0.485 ;
        RECT 1.26 0.215 1.4 0.305 ;
      LAYER MET2 ;
        RECT 5.05 0.23 5.15 0.76 ;
      LAYER VIA1 ;
        RECT 5.055 0.455 5.145 0.545 ;
    END
  END Z
  OBS
    LAYER MET1 ;
      RECT 3.29 1.065 5.38 1.155 ;
      RECT 3.29 0.9 3.38 1.155 ;
      RECT 1.26 0.9 3.38 0.99 ;
      RECT 0.755 1.06 0.9 1.15 ;
      RECT 0.755 0.85 0.845 1.15 ;
      RECT 0.26 0.85 0.845 0.94 ;
      RECT 0.285 0.33 0.375 0.94 ;
      RECT 1.115 0.64 2.93 0.73 ;
      RECT 1.115 0.395 1.205 0.73 ;
      RECT 0.285 0.395 1.205 0.485 ;
  END
END NOR2BX16H7R

MACRO NOR2BX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BX1H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.32 0.975 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.81 -0.08 0.95 0.175 ;
        RECT 0.295 -0.08 0.435 0.335 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.345 0.855 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.55 0.775 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.755 0.885 0.955 0.975 ;
        RECT 0.865 0.265 0.955 0.975 ;
        RECT 0.855 0.825 0.955 0.975 ;
        RECT 0.545 0.265 0.955 0.355 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Z
  OBS
    LAYER MET1 ;
      RECT 0.045 0.945 0.185 1.035 ;
      RECT 0.045 0.26 0.135 1.035 ;
      RECT 0.455 0.445 0.545 0.645 ;
      RECT 0.045 0.445 0.545 0.535 ;
      RECT 0.045 0.26 0.185 0.35 ;
  END
END NOR2BX1H7R

MACRO NOR2BX1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BX1P4H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.32 1.019 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.815 -0.08 0.955 0.33 ;
        RECT 0.32 -0.08 0.41 0.34 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.345 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.635 0.6 0.775 0.795 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.885 0.955 1.175 ;
        RECT 0.865 0.42 0.955 1.175 ;
        RECT 0.635 0.42 0.955 0.51 ;
        RECT 0.755 0.885 0.955 0.975 ;
        RECT 0.635 0.265 0.725 0.51 ;
        RECT 0.545 0.265 0.725 0.355 ;
      LAYER MET2 ;
        RECT 0.85 0.84 0.95 1.22 ;
      LAYER VIA1 ;
        RECT 0.855 1.055 0.945 1.145 ;
    END
  END Z
  OBS
    LAYER MET1 ;
      RECT 0.045 0.989 0.185 1.079 ;
      RECT 0.045 0.24 0.135 1.079 ;
      RECT 0.455 0.445 0.545 0.66 ;
      RECT 0.045 0.445 0.545 0.535 ;
      RECT 0.045 0.24 0.185 0.33 ;
  END
END NOR2BX1P4H7R

MACRO NOR2BX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BX2H7R 0 0 ;
  SIZE 1.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.2 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.2 0.08 ;
        RECT 0.835 -0.08 0.925 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.345 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.615 0.775 0.84 ;
      LAYER MET2 ;
        RECT 0.65 0.6 0.75 1.135 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.865 0.435 0.955 0.965 ;
        RECT 0.655 0.435 0.955 0.525 ;
        RECT 0.655 0.225 0.745 0.525 ;
        RECT 0.545 0.225 0.745 0.315 ;
      LAYER MET2 ;
        RECT 0.65 0.18 0.75 0.385 ;
      LAYER VIA1 ;
        RECT 0.655 0.255 0.745 0.345 ;
    END
  END Z
  OBS
    LAYER MET1 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 0.455 0.445 0.545 0.755 ;
      RECT 0.045 0.445 0.545 0.535 ;
      RECT 0.045 0.23 0.185 0.32 ;
  END
END NOR2BX2H7R

MACRO NOR2BX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BX3H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 0.795 1.08 0.935 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.565 -0.08 1.655 0.345 ;
        RECT 1.065 -0.08 1.155 0.345 ;
        RECT 0.82 -0.08 0.91 0.345 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.36 0.825 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.635 1.225 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.315 0.295 1.405 1.045 ;
        RECT 0.64 0.455 1.405 0.545 ;
        RECT 0.64 0.24 0.73 0.545 ;
        RECT 0.545 0.24 0.73 0.33 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END Z
  OBS
    LAYER MET1 ;
      RECT 1.065 1.135 1.655 1.225 ;
      RECT 1.565 1.055 1.655 1.225 ;
      RECT 1.065 0.9 1.155 1.225 ;
      RECT 0.57 0.9 0.66 1.045 ;
      RECT 0.57 0.9 1.155 0.99 ;
      RECT 0.045 0.96 0.185 1.05 ;
      RECT 0.045 0.29 0.135 1.05 ;
      RECT 0.46 0.64 0.815 0.73 ;
      RECT 0.46 0.42 0.55 0.73 ;
      RECT 0.045 0.42 0.55 0.51 ;
      RECT 0.045 0.29 0.185 0.51 ;
  END
END NOR2BX3H7R

MACRO NOR2BX4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BX4H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 0.97 1.08 1.11 1.48 ;
        RECT 0.495 1.07 0.585 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.74 -0.08 1.83 0.345 ;
        RECT 1.24 -0.08 1.33 0.345 ;
        RECT 0.995 -0.08 1.085 0.345 ;
        RECT 0.495 -0.08 0.585 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.395 0.6 0.545 0.78 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.22 0.635 1.4 0.785 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.49 0.37 1.58 0.95 ;
        RECT 0.815 0.455 1.58 0.545 ;
        RECT 0.815 0.24 0.905 0.545 ;
        RECT 0.72 0.24 0.905 0.33 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END Z
  OBS
    LAYER MET1 ;
      RECT 1.265 1.04 1.855 1.13 ;
      RECT 1.265 0.9 1.355 1.13 ;
      RECT 0.72 0.9 1.355 0.99 ;
      RECT 0.215 1.04 0.36 1.13 ;
      RECT 0.215 0.33 0.305 1.13 ;
      RECT 0.635 0.64 0.99 0.73 ;
      RECT 0.635 0.42 0.725 0.73 ;
      RECT 0.215 0.42 0.725 0.51 ;
      RECT 0.215 0.33 0.36 0.51 ;
  END
END NOR2BX4H7R

MACRO NOR2BX6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BX6H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 1.032 1.07 1.122 1.48 ;
        RECT 0.532 1.07 0.622 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 2.007 -0.08 2.147 0.32 ;
        RECT 1.532 -0.08 1.622 0.33 ;
        RECT 1.032 -0.08 1.122 0.33 ;
        RECT 0.532 -0.08 0.622 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.437 0.6 0.572 0.8 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.425 0.655 1.965 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.507 0.885 2.147 0.975 ;
        RECT 2.055 0.42 2.147 0.975 ;
        RECT 0.852 0.42 2.147 0.51 ;
        RECT 1.782 0.37 1.872 0.51 ;
        RECT 1.282 0.37 1.372 0.51 ;
        RECT 0.852 0.24 0.942 0.51 ;
        RECT 0.757 0.24 0.942 0.33 ;
      LAYER MET2 ;
        RECT 2.05 0.23 2.15 0.76 ;
      LAYER VIA1 ;
        RECT 2.055 0.455 2.145 0.545 ;
    END
  END Z
  OBS
    LAYER MET1 ;
      RECT 1.302 1.065 1.897 1.155 ;
      RECT 1.302 0.89 1.397 1.155 ;
      RECT 0.757 0.89 1.397 0.98 ;
      RECT 0.257 0.89 0.397 0.98 ;
      RECT 0.257 0.33 0.347 0.98 ;
      RECT 0.672 0.64 1.027 0.73 ;
      RECT 0.672 0.42 0.762 0.73 ;
      RECT 0.257 0.42 0.762 0.51 ;
      RECT 0.257 0.33 0.397 0.51 ;
  END
END NOR2BX6H7R

MACRO NOR2BX8H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BX8H7R 0 0 ;
  SIZE 3.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.2 1.48 ;
        RECT 1.545 1.08 1.685 1.48 ;
        RECT 1.07 1.07 1.16 1.48 ;
        RECT 0.57 1.07 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.2 0.08 ;
        RECT 2.81 -0.08 2.95 0.305 ;
        RECT 2.302 -0.08 2.442 0.305 ;
        RECT 1.79 -0.08 1.93 0.305 ;
        RECT 1.045 -0.08 1.185 0.305 ;
        RECT 0.57 -0.08 0.66 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.615 0.59 0.815 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.025 0.655 2.765 0.745 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END B
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.06 0.885 2.945 0.975 ;
        RECT 2.855 0.395 2.945 0.975 ;
        RECT 0.86 0.395 2.945 0.485 ;
        RECT 0.86 0.24 0.95 0.485 ;
        RECT 0.795 0.24 0.95 0.33 ;
      LAYER MET2 ;
        RECT 2.85 0.23 2.95 0.76 ;
      LAYER VIA1 ;
        RECT 2.855 0.455 2.945 0.545 ;
    END
  END Z
  OBS
    LAYER MET1 ;
      RECT 1.86 1.065 2.95 1.155 ;
      RECT 1.86 0.89 1.95 1.155 ;
      RECT 0.795 0.89 1.95 0.98 ;
      RECT 0.275 0.905 0.435 0.995 ;
      RECT 0.275 0.33 0.365 0.995 ;
      RECT 0.68 0.64 1.465 0.73 ;
      RECT 0.68 0.435 0.77 0.73 ;
      RECT 0.275 0.435 0.77 0.525 ;
      RECT 0.275 0.33 0.435 0.525 ;
  END
END NOR2BX8H7R

MACRO NOR2X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X0P5H7R 0 0 ;
  SIZE 0.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.8 1.48 ;
        RECT 0.07 0.865 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.8 0.08 ;
        RECT 0.615 -0.08 0.755 0.175 ;
        RECT 0.07 -0.08 0.16 0.38 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.18 0.61 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.64 0.545 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.64 0.275 0.745 0.99 ;
        RECT 0.345 0.275 0.745 0.365 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END Y
END NOR2X0P5H7R

MACRO NOR2X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X0P7H7R 0 0 ;
  SIZE 0.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.8 1.48 ;
        RECT 0.07 0.897 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.8 0.08 ;
        RECT 0.615 -0.08 0.755 0.21 ;
        RECT 0.07 -0.08 0.16 0.38 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.365 0.625 0.545 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.64 0.3 0.745 0.975 ;
        RECT 0.345 0.3 0.745 0.39 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END Y
END NOR2X0P7H7R

MACRO NOR2X12H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X12H7R 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.8 1.48 ;
        RECT 1.547 1.095 1.687 1.48 ;
        RECT 1.047 1.095 1.187 1.48 ;
        RECT 0.547 1.095 0.687 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.8 0.08 ;
        RECT 3.297 -0.08 3.437 0.305 ;
        RECT 2.797 -0.08 2.937 0.305 ;
        RECT 2.297 -0.08 2.437 0.305 ;
        RECT 1.797 -0.08 1.937 0.305 ;
        RECT 1.297 -0.08 1.437 0.305 ;
        RECT 0.797 -0.08 0.937 0.305 ;
        RECT 0.322 -0.08 0.412 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.617 0.655 1.757 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.977 0.655 3.117 0.745 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.047 0.885 3.345 0.975 ;
        RECT 3.255 0.395 3.345 0.975 ;
        RECT 0.547 0.395 3.345 0.485 ;
      LAYER MET2 ;
        RECT 3.25 0.23 3.35 0.76 ;
      LAYER VIA1 ;
        RECT 3.255 0.455 3.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.822 1.07 3.437 1.16 ;
      RECT 1.822 0.915 1.912 1.16 ;
      RECT 0.297 0.915 1.912 1.005 ;
  END
END NOR2X12H7R

MACRO NOR2X16H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X16H7R 0 0 ;
  SIZE 4.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.8 1.48 ;
        RECT 2.047 1.095 2.187 1.48 ;
        RECT 1.547 1.095 1.687 1.48 ;
        RECT 1.047 1.095 1.187 1.48 ;
        RECT 0.547 1.095 0.687 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.8 0.08 ;
        RECT 4.297 -0.08 4.437 0.305 ;
        RECT 3.797 -0.08 3.937 0.305 ;
        RECT 3.297 -0.08 3.437 0.305 ;
        RECT 2.797 -0.08 2.937 0.305 ;
        RECT 2.297 -0.08 2.437 0.305 ;
        RECT 1.797 -0.08 1.937 0.305 ;
        RECT 1.297 -0.08 1.437 0.305 ;
        RECT 0.797 -0.08 0.937 0.305 ;
        RECT 0.322 -0.08 0.412 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.517 0.655 2.257 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.477 0.655 4.017 0.745 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.547 0.885 4.345 0.975 ;
        RECT 4.255 0.395 4.345 0.975 ;
        RECT 0.547 0.395 4.345 0.485 ;
      LAYER MET2 ;
        RECT 4.25 0.425 4.35 0.96 ;
      LAYER VIA1 ;
        RECT 4.255 0.655 4.345 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.322 1.065 4.437 1.155 ;
      RECT 2.322 0.915 2.412 1.155 ;
      RECT 0.297 0.915 2.412 1.005 ;
  END
END NOR2X16H7R

MACRO NOR2X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X1H7R 0 0 ;
  SIZE 0.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.8 1.48 ;
        RECT 0.07 0.89 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.8 0.08 ;
        RECT 0.635 -0.08 0.725 0.21 ;
        RECT 0.07 -0.08 0.16 0.39 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.58 0.545 0.84 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.595 0.935 0.745 1.025 ;
        RECT 0.655 0.35 0.745 1.025 ;
        RECT 0.305 0.35 0.745 0.44 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END Y
END NOR2X1H7R

MACRO NOR2X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X1P4H7R 0 0 ;
  SIZE 0.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.8 1.48 ;
        RECT 0.07 1.004 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.8 0.08 ;
        RECT 0.635 -0.08 0.725 0.26 ;
        RECT 0.07 -0.08 0.16 0.355 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.58 0.545 0.78 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.545 0.935 0.745 1.025 ;
        RECT 0.655 0.35 0.745 1.025 ;
        RECT 0.295 0.35 0.745 0.44 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END Y
END NOR2X1P4H7R

MACRO NOR2X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X2H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.31 1.215 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.15 -0.08 1.24 0.43 ;
        RECT 0.59 -0.08 0.73 0.175 ;
        RECT 0.07 -0.08 0.16 0.43 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.195 0.655 0.535 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.55 1.345 0.775 ;
        RECT 0.945 0.55 1.345 0.64 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.75 0.995 1.04 ;
        RECT 0.3 0.315 0.995 0.405 ;
        RECT 0.655 0.75 0.995 0.84 ;
        RECT 0.655 0.315 0.745 0.84 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.6 1.135 1.24 1.225 ;
      RECT 1.15 0.98 1.24 1.225 ;
      RECT 0.6 0.965 0.69 1.225 ;
      RECT 0.045 0.965 0.69 1.055 ;
  END
END NOR2X2H7R

MACRO NOR2X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X3H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.31 1.175 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.15 -0.08 1.24 0.375 ;
        RECT 0.59 -0.08 0.73 0.26 ;
        RECT 0.07 -0.08 0.16 0.375 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.195 0.655 0.535 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.605 1.145 0.795 ;
        RECT 0.945 0.605 1.145 0.695 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.3 0.35 0.995 0.44 ;
        RECT 0.765 0.855 0.975 0.945 ;
        RECT 0.765 0.35 0.855 0.945 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.6 1.065 1.24 1.155 ;
      RECT 1.15 0.98 1.24 1.155 ;
      RECT 0.045 0.995 0.69 1.085 ;
  END
END NOR2X3H7R

MACRO NOR2X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X4H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 0.87 1.155 1.01 1.48 ;
        RECT 0.31 1.155 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 2.22 -0.08 2.31 0.435 ;
        RECT 1.68 -0.08 1.82 0.175 ;
        RECT 1.15 -0.08 1.29 0.175 ;
        RECT 0.59 -0.08 0.73 0.175 ;
        RECT 0.07 -0.08 0.16 0.43 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.195 0.635 1.135 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.255 0.535 2.345 0.775 ;
        RECT 1.635 0.535 2.345 0.625 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.31 0.315 2.085 0.405 ;
        RECT 1.915 0.745 2.055 1.04 ;
        RECT 1.415 0.745 2.055 0.835 ;
        RECT 1.415 0.745 1.561 1.04 ;
        RECT 1.415 0.315 1.545 1.04 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.16 1.135 2.31 1.225 ;
      RECT 2.22 0.961 2.31 1.225 ;
      RECT 1.69 0.94 1.78 1.225 ;
      RECT 1.16 0.965 1.25 1.225 ;
      RECT 0.045 0.965 1.25 1.055 ;
  END
END NOR2X4H7R

MACRO NOR2X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X6H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 0.87 1.2 1.01 1.48 ;
        RECT 0.31 1.2 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 2.22 -0.08 2.31 0.375 ;
        RECT 1.68 -0.08 1.82 0.26 ;
        RECT 1.15 -0.08 1.29 0.26 ;
        RECT 0.59 -0.08 0.73 0.26 ;
        RECT 0.07 -0.08 0.16 0.375 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.655 0.965 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.395 0.655 2.135 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.325 0.35 2.114 0.44 ;
        RECT 1.945 0.84 2.085 0.975 ;
        RECT 1.055 0.84 2.085 0.93 ;
        RECT 1.415 0.84 1.555 0.975 ;
        RECT 1.055 0.35 1.145 0.93 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.185 1.065 2.31 1.155 ;
      RECT 2.22 0.98 2.31 1.155 ;
      RECT 0.07 1.02 1.275 1.11 ;
      RECT 1.665 1.02 1.805 1.155 ;
      RECT 0.07 0.97 0.16 1.11 ;
  END
END NOR2X6H7R

MACRO NOR2X8H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X8H7R 0 0 ;
  SIZE 2.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.8 1.48 ;
        RECT 1.072 1.07 1.162 1.48 ;
        RECT 0.572 1.07 0.662 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.8 0.08 ;
        RECT 2.297 -0.08 2.437 0.305 ;
        RECT 1.797 -0.08 1.937 0.305 ;
        RECT 1.297 -0.08 1.437 0.305 ;
        RECT 0.797 -0.08 0.937 0.305 ;
        RECT 0.322 -0.08 0.412 0.375 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.517 0.655 1.257 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.48 0.655 2.02 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.547 0.885 2.345 0.975 ;
        RECT 2.255 0.395 2.345 0.975 ;
        RECT 0.572 0.395 2.345 0.485 ;
        RECT 0.572 0.345 0.662 0.485 ;
      LAYER MET2 ;
        RECT 2.25 0.23 2.35 0.76 ;
      LAYER VIA1 ;
        RECT 2.255 0.455 2.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.322 1.065 2.437 1.155 ;
      RECT 1.322 0.89 1.412 1.155 ;
      RECT 0.297 0.89 1.412 0.98 ;
  END
END NOR2X8H7R

MACRO NOR3BX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BX0P5H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.32 0.88 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.885 -0.08 1.025 0.345 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.575 0.385 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.625 0.835 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.625 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.135 0.865 1.345 0.955 ;
        RECT 1.255 0.425 1.345 0.955 ;
        RECT 0.66 0.435 1.345 0.525 ;
        RECT 1.16 0.425 1.345 0.525 ;
        RECT 1.16 0.245 1.25 0.525 ;
        RECT 0.66 0.26 0.75 0.525 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.27 0.16 0.965 ;
      RECT 0.48 0.27 0.57 0.595 ;
      RECT 0.045 0.27 0.57 0.36 ;
  END
END NOR3BX0P5H7R

MACRO NOR3BX0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BX0P7H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.395 0.97 0.485 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.935 -0.08 1.075 0.345 ;
        RECT 0.335 -0.08 0.475 0.18 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.575 0.385 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.765 0.625 0.945 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.673 1.145 0.975 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.24 0.225 1.345 1.023 ;
        RECT 0.695 0.435 1.345 0.525 ;
        RECT 0.695 0.285 0.785 0.525 ;
      LAYER MET2 ;
        RECT 1.25 0.18 1.35 0.56 ;
      LAYER VIA1 ;
        RECT 1.255 0.255 1.345 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.27 0.16 1.055 ;
      RECT 0.51 0.27 0.6 0.62 ;
      RECT 0.045 0.27 0.6 0.36 ;
  END
END NOR3BX0P7H7R

MACRO NOR3BX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BX1H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.425 0.877 0.565 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.95 -0.08 1.09 0.175 ;
        RECT 0.42 -0.08 0.56 0.175 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.515 0.36 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.81 0.575 0.945 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.63 1.145 0.975 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.24 0.295 1.345 1.037 ;
        RECT 0.685 0.295 1.345 0.385 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.075 0.878 0.28 0.968 ;
      RECT 0.075 0.275 0.165 0.968 ;
      RECT 0.505 0.275 0.595 0.66 ;
      RECT 0.075 0.275 0.595 0.365 ;
  END
END NOR3BX1H7R

MACRO NOR3BX1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BX1P4H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.395 0.97 0.485 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.935 -0.08 1.075 0.305 ;
        RECT 0.36 -0.08 0.45 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.625 0.4 0.805 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.795 0.595 0.945 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.581 1.145 0.975 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.24 0.3 1.345 0.931 ;
        RECT 0.695 0.401 1.345 0.491 ;
        RECT 0.695 0.315 0.785 0.491 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.205 0.16 1.055 ;
      RECT 0.51 0.445 0.6 0.65 ;
      RECT 0.07 0.445 0.6 0.535 ;
  END
END NOR3BX1P4H7R

MACRO NOR3BX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BX2H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 0.45 0.85 0.74 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 2.02 -0.08 2.11 0.39 ;
        RECT 1.505 -0.08 1.595 0.2 ;
        RECT 0.975 -0.08 1.065 0.2 ;
        RECT 0.42 -0.08 0.56 0.175 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.55 0.375 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.085 0.645 1.425 0.745 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.425 0.855 1.675 0.945 ;
        RECT 1.585 0.595 1.675 0.945 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.77 0.805 2.06 1.145 ;
        RECT 1.77 0.29 1.885 1.145 ;
        RECT 0.685 0.29 1.885 0.38 ;
      LAYER MET2 ;
        RECT 1.85 0.625 1.95 1.16 ;
      LAYER VIA1 ;
        RECT 1.855 0.855 1.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.075 0.87 0.28 0.96 ;
      RECT 0.075 0.275 0.165 0.96 ;
      RECT 0.505 0.545 0.925 0.635 ;
      RECT 0.505 0.275 0.595 0.635 ;
      RECT 0.075 0.275 0.595 0.365 ;
  END
END NOR3BX2H7R

MACRO NOR3BX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BX3H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 0.92 1.035 1.01 1.48 ;
        RECT 0.42 1.05 0.51 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 2.15 -0.08 2.24 0.375 ;
        RECT 1.55 -0.08 1.69 0.26 ;
        RECT 0.95 -0.08 1.09 0.26 ;
        RECT 0.42 -0.08 0.56 0.23 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.55 0.375 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.195 0.655 1.535 0.745 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.625 0.655 1.895 0.755 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.9 0.855 2.145 0.945 ;
        RECT 2.055 0.494 2.145 0.945 ;
        RECT 1.979 0.449 2.101 0.501 ;
        RECT 1.941 0.411 2.055 0.459 ;
        RECT 2.025 0.494 2.145 0.539 ;
        RECT 0.685 0.373 2.025 0.44 ;
        RECT 1.9 0.855 1.99 1.025 ;
        RECT 0.685 0.35 1.979 0.44 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.15 1.14 2.24 1.23 ;
      RECT 2.15 1.035 2.24 1.23 ;
      RECT 1.65 1.05 1.74 1.23 ;
      RECT 1.15 1.035 1.24 1.23 ;
      RECT 1.4 0.855 1.49 1.025 ;
      RECT 0.67 0.855 0.76 1.025 ;
      RECT 0.67 0.855 1.49 0.945 ;
      RECT 0.075 0.94 0.28 1.03 ;
      RECT 0.075 0.32 0.165 1.03 ;
      RECT 0.505 0.58 0.875 0.67 ;
      RECT 0.505 0.32 0.595 0.67 ;
      RECT 0.075 0.32 0.595 0.41 ;
  END
END NOR3BX3H7R

MACRO NOR3BX4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BX4H7R 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.8 1.48 ;
        RECT 1.095 1.005 1.235 1.48 ;
        RECT 0.6 0.98 0.69 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.8 0.08 ;
        RECT 3.25 -0.08 3.39 0.175 ;
        RECT 2.715 -0.08 2.855 0.175 ;
        RECT 2.2 -0.08 2.34 0.175 ;
        RECT 1.665 -0.08 1.805 0.175 ;
        RECT 1.15 -0.08 1.29 0.175 ;
        RECT 0.63 -0.08 0.72 0.35 ;
        RECT 0.385 -0.08 0.475 0.35 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.315 0.62 0.545 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.85 0.52 2.39 0.61 ;
        RECT 2.225 0.455 2.39 0.61 ;
      LAYER MET2 ;
        RECT 2.25 0.23 2.35 0.76 ;
      LAYER VIA1 ;
        RECT 2.255 0.455 2.345 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.825 0.52 3.37 0.61 ;
        RECT 2.825 0.455 2.975 0.61 ;
      LAYER MET2 ;
        RECT 2.85 0.23 2.95 0.76 ;
      LAYER VIA1 ;
        RECT 2.855 0.455 2.945 0.545 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.54 0.225 3.745 0.375 ;
        RECT 3.51 0.825 3.63 1.1 ;
        RECT 3.54 0.225 3.63 1.1 ;
        RECT 0.885 0.265 3.745 0.355 ;
        RECT 2.985 0.825 3.63 0.915 ;
      LAYER MET2 ;
        RECT 3.65 0.18 3.75 0.56 ;
      LAYER VIA1 ;
        RECT 3.655 0.255 3.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.92 1.005 3.375 1.095 ;
      RECT 2.445 0.81 2.535 1.095 ;
      RECT 1.37 0.825 1.46 1.1 ;
      RECT 0.845 0.825 2.31 0.915 ;
      RECT 0.135 0.31 0.225 0.945 ;
      RECT 0.705 0.515 1.315 0.605 ;
      RECT 0.135 0.44 0.795 0.53 ;
  END
END NOR3BX4H7R

MACRO NOR3BX6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BX6H7R 0 0 ;
  SIZE 3.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.4 1.48 ;
        RECT 1.035 1.07 1.125 1.48 ;
        RECT 0.535 1.07 0.625 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.4 0.08 ;
        RECT 3.025 -0.08 3.115 0.345 ;
        RECT 2.525 -0.08 2.615 0.33 ;
        RECT 2.025 -0.08 2.115 0.33 ;
        RECT 1.525 -0.08 1.615 0.345 ;
        RECT 1.035 -0.08 1.125 0.33 ;
        RECT 0.535 -0.08 0.625 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.435 0.6 0.585 0.78 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.67 0.655 2.21 0.745 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.42 0.655 2.96 0.745 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.5 1.065 3.145 1.155 ;
        RECT 3.055 0.455 3.145 1.155 ;
        RECT 0.855 0.455 3.145 0.545 ;
        RECT 2.775 0.37 2.865 0.545 ;
        RECT 2.275 0.37 2.365 0.545 ;
        RECT 1.775 0.37 1.865 0.545 ;
        RECT 1.285 0.355 1.375 0.545 ;
        RECT 0.855 0.24 0.945 0.545 ;
        RECT 0.76 0.24 0.945 0.33 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.55 1.065 2.14 1.155 ;
      RECT 1.55 0.89 1.64 1.155 ;
      RECT 0.76 0.89 1.64 0.98 ;
      RECT 0.255 0.865 0.4 0.955 ;
      RECT 0.255 0.33 0.345 0.955 ;
      RECT 0.675 0.64 1.23 0.73 ;
      RECT 0.675 0.42 0.765 0.73 ;
      RECT 0.255 0.42 0.765 0.51 ;
      RECT 0.255 0.33 0.4 0.51 ;
      RECT 1.75 0.885 2.89 0.975 ;
  END
END NOR3BX6H7R

MACRO NOR3X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X0P5H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.045 0.91 0.185 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.545 -0.08 0.685 0.305 ;
        RECT 0.045 -0.08 0.185 0.32 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.42 0.635 0.545 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.635 0.575 0.76 0.815 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.82 0.885 0.945 1.03 ;
        RECT 0.85 0.395 0.945 1.03 ;
        RECT 0.82 0.205 0.915 0.485 ;
        RECT 0.32 0.395 0.945 0.485 ;
        RECT 0.32 0.205 0.41 0.485 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END Y
END NOR3X0P5H7R

MACRO NOR3X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X0P7H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.07 0.917 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.545 -0.08 0.685 0.305 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.625 0.545 0.825 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.635 0.745 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.835 0.225 0.945 0.985 ;
        RECT 0.32 0.395 0.945 0.485 ;
        RECT 0.32 0.245 0.41 0.485 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.56 ;
      LAYER VIA1 ;
        RECT 0.855 0.255 0.945 0.345 ;
    END
  END Y
END NOR3X0P7H7R

MACRO NOR3X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X1H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.07 0.91 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.565 -0.08 0.705 0.345 ;
        RECT 0.075 -0.08 0.165 0.42 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.63 0.545 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.615 0.765 0.865 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.84 0.96 0.945 1.1 ;
        RECT 0.855 0.305 0.945 1.1 ;
        RECT 0.33 0.435 0.945 0.525 ;
        RECT 0.84 0.305 0.945 0.525 ;
        RECT 0.33 0.29 0.42 0.525 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END Y
END NOR3X1H7R

MACRO NOR3X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X1P4H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.545 -0.08 0.685 0.305 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.625 0.545 0.825 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.641 0.745 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.835 0.3 0.945 1.031 ;
        RECT 0.32 0.395 0.945 0.485 ;
        RECT 0.32 0.315 0.41 0.485 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END Y
END NOR3X1P4H7R

MACRO NOR3X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X2H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 0.07 0.855 0.36 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.64 -0.08 1.73 0.365 ;
        RECT 1.1 -0.08 1.24 0.175 ;
        RECT 0.57 -0.08 0.71 0.175 ;
        RECT 0.075 -0.08 0.165 0.365 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.175 0.65 0.515 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.705 0.655 1.045 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.245 0.615 1.365 0.84 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.265 1.545 1.165 ;
        RECT 0.305 0.265 1.545 0.355 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END Y
END NOR3X2H7R

MACRO NOR3X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X3H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.64 -0.08 1.73 0.365 ;
        RECT 1.1 -0.08 1.24 0.25 ;
        RECT 0.57 -0.08 0.71 0.25 ;
        RECT 0.075 -0.08 0.165 0.365 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.175 0.655 0.515 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.705 0.655 1.045 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.295 0.655 1.635 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.8 0.455 1.89 1.06 ;
        RECT 1.275 0.915 1.89 1.005 ;
        RECT 1.455 0.455 1.89 0.545 ;
        RECT 1.455 0.34 1.545 0.545 ;
        RECT 0.305 0.34 1.545 0.43 ;
        RECT 1.275 0.915 1.415 1.035 ;
      LAYER MET2 ;
        RECT 1.65 0.23 1.75 0.76 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.795 1.125 1.665 1.215 ;
      RECT 1.525 1.095 1.665 1.215 ;
      RECT 0.795 1.095 0.935 1.215 ;
      RECT 0.07 0.915 0.16 1.06 ;
      RECT 0.57 0.915 0.66 1.045 ;
      RECT 1.045 0.915 1.185 1.035 ;
      RECT 0.07 0.915 1.185 1.005 ;
  END
END NOR3X3H7R

MACRO NOR3X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X4H7R 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.8 1.48 ;
        RECT 1.09 1.225 1.23 1.48 ;
        RECT 0.56 1.225 0.7 1.48 ;
        RECT 0.07 0.93 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.8 0.08 ;
        RECT 3.45 -0.08 3.54 0.415 ;
        RECT 2.91 -0.08 3.05 0.175 ;
        RECT 2.38 -0.08 2.52 0.175 ;
        RECT 1.85 -0.08 1.99 0.175 ;
        RECT 1.32 -0.08 1.46 0.175 ;
        RECT 1.09 -0.08 1.23 0.175 ;
        RECT 0.56 -0.08 0.7 0.175 ;
        RECT 0.07 -0.08 0.16 0.415 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.655 0.965 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.55 0.655 2.29 0.745 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.695 0.655 3.235 0.745 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.515 0.855 3.315 0.985 ;
        RECT 0.295 0.3 3.315 0.39 ;
        RECT 2.515 0.3 2.605 0.985 ;
      LAYER MET2 ;
        RECT 2.65 0.63 2.75 1.16 ;
      LAYER VIA1 ;
        RECT 2.655 0.855 2.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.32 1.11 3.54 1.2 ;
      RECT 3.45 0.905 3.54 1.2 ;
      RECT 0.295 0.93 2.255 1.02 ;
  END
END NOR3X4H7R

MACRO NOR3X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X6H7R 0 0 ;
  SIZE 3 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3 1.48 ;
        RECT 0.825 1.07 0.915 1.48 ;
        RECT 0.325 1.055 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3 0.08 ;
        RECT 2.3 -0.08 2.44 0.305 ;
        RECT 1.8 -0.08 1.94 0.305 ;
        RECT 1.3 -0.08 1.44 0.305 ;
        RECT 0.8 -0.08 0.94 0.305 ;
        RECT 0.325 -0.08 0.415 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.47 0.655 1.01 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.23 0.655 1.77 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.97 0.655 2.51 0.745 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.05 0.885 2.745 0.975 ;
        RECT 2.655 0.395 2.745 0.975 ;
        RECT 2.575 0.205 2.665 0.485 ;
        RECT 0.55 0.395 2.745 0.485 ;
      LAYER MET2 ;
        RECT 2.65 0.23 2.75 0.76 ;
      LAYER VIA1 ;
        RECT 2.655 0.455 2.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.3 1.08 2.44 1.17 ;
      RECT 0.55 0.885 1.69 0.975 ;
  END
END NOR3X6H7R

MACRO NOR3X8H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X8H7R 0 0 ;
  SIZE 4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4 1.48 ;
        RECT 1.075 1.07 1.165 1.48 ;
        RECT 0.575 1.07 0.665 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4 0.08 ;
        RECT 3.31 -0.08 3.45 0.305 ;
        RECT 2.81 -0.08 2.95 0.305 ;
        RECT 2.3 -0.08 2.44 0.305 ;
        RECT 1.8 -0.08 1.94 0.305 ;
        RECT 1.3 -0.08 1.44 0.305 ;
        RECT 0.8 -0.08 0.94 0.305 ;
        RECT 0.325 -0.08 0.415 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.495 0.655 1.235 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.48 0.655 2.22 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.745 0.655 3.485 0.745 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.81 0.885 3.745 0.975 ;
        RECT 3.655 0.395 3.745 0.975 ;
        RECT 3.585 0.205 3.675 0.485 ;
        RECT 0.55 0.395 3.745 0.485 ;
      LAYER MET2 ;
        RECT 3.65 0.23 3.75 0.76 ;
      LAYER VIA1 ;
        RECT 3.655 0.455 3.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.55 1.08 3.7 1.17 ;
      RECT 0.3 0.885 2.44 0.975 ;
  END
END NOR3X8H7R

MACRO NOR4BBX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BBX0P5H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.835 0.975 1.925 1.48 ;
        RECT 0.325 0.99 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.355 -0.08 1.445 0.37 ;
        RECT 0.815 -0.08 0.955 0.175 ;
        RECT 0.325 -0.08 0.415 0.365 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.655 0.375 0.835 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.815 0.615 1.95 0.815 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.815 0.445 1.04 0.565 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.365 0.625 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.13 0.96 1.47 1.05 ;
        RECT 1.13 0.255 1.22 1.05 ;
        RECT 0.55 0.265 1.22 0.355 ;
        RECT 1.025 0.255 1.22 0.355 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.56 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.675 1.14 1.675 1.23 ;
      RECT 1.585 0.878 1.675 1.23 ;
      RECT 1.631 0.853 1.675 1.23 ;
      RECT 0.675 0.725 0.765 1.23 ;
      RECT 1.585 0.878 1.721 0.916 ;
      RECT 1.635 0.265 1.725 0.891 ;
      RECT 1.635 0.265 1.95 0.355 ;
      RECT 0.045 0.96 0.19 1.05 ;
      RECT 0.045 0.265 0.135 1.05 ;
      RECT 0.045 0.475 0.565 0.565 ;
      RECT 0.045 0.265 0.14 0.565 ;
      RECT 0.045 0.265 0.19 0.355 ;
  END
END NOR4BBX0P5H7R

MACRO NOR4BBX0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BBX0P7H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.835 0.975 1.925 1.48 ;
        RECT 0.325 0.99 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.355 -0.08 1.445 0.37 ;
        RECT 0.815 -0.08 0.955 0.175 ;
        RECT 0.3 -0.08 0.44 0.34 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.345 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.815 0.615 1.95 0.815 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.455 1.025 0.595 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.365 0.625 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.13 0.928 1.47 1.018 ;
        RECT 1.13 0.255 1.22 1.018 ;
        RECT 0.55 0.265 1.22 0.355 ;
        RECT 1.025 0.255 1.22 0.355 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.56 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.675 1.108 1.675 1.198 ;
      RECT 1.585 0.878 1.675 1.198 ;
      RECT 1.631 0.853 1.675 1.198 ;
      RECT 0.675 0.693 0.765 1.198 ;
      RECT 1.585 0.878 1.721 0.916 ;
      RECT 1.635 0.265 1.725 0.891 ;
      RECT 1.635 0.265 1.95 0.355 ;
      RECT 0.045 0.96 0.19 1.05 ;
      RECT 0.045 0.265 0.135 1.05 ;
      RECT 0.45 0.445 0.54 0.615 ;
      RECT 0.045 0.445 0.54 0.535 ;
      RECT 0.045 0.265 0.14 0.535 ;
      RECT 0.045 0.265 0.19 0.355 ;
  END
END NOR4BBX0P7H7R

MACRO NOR4BBX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BBX1H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.835 0.975 1.925 1.48 ;
        RECT 0.325 0.99 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.39 -0.08 1.48 0.365 ;
        RECT 0.815 -0.08 0.955 0.175 ;
        RECT 0.3 -0.08 0.44 0.34 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.345 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.815 0.6 1.95 0.8 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.955 0.455 1.045 0.65 ;
        RECT 0.825 0.455 1.045 0.545 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.365 0.625 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.155 0.88 1.47 0.97 ;
        RECT 1.155 0.255 1.245 0.97 ;
        RECT 0.55 0.265 1.245 0.355 ;
        RECT 1.025 0.255 1.245 0.355 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.56 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.715 1.06 1.675 1.15 ;
      RECT 1.585 0.863 1.675 1.15 ;
      RECT 1.631 0.838 1.675 1.15 ;
      RECT 0.715 0.645 0.805 1.15 ;
      RECT 1.585 0.863 1.721 0.901 ;
      RECT 1.635 0.265 1.725 0.876 ;
      RECT 1.635 0.265 1.95 0.355 ;
      RECT 0.045 0.96 0.19 1.05 ;
      RECT 0.045 0.265 0.135 1.05 ;
      RECT 0.455 0.445 0.545 0.65 ;
      RECT 0.045 0.445 0.545 0.535 ;
      RECT 0.045 0.265 0.14 0.535 ;
      RECT 0.045 0.265 0.19 0.355 ;
  END
END NOR4BBX1H7R

MACRO NOR4BBX1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BBX1P4H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.835 0.975 1.925 1.48 ;
        RECT 0.325 1.055 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.39 -0.08 1.48 0.33 ;
        RECT 0.84 -0.08 0.93 0.33 ;
        RECT 0.325 -0.08 0.415 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.345 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.815 0.6 1.95 0.8 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.855 1.035 0.945 ;
        RECT 0.945 0.706 1.035 0.945 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.365 0.625 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.125 0.916 1.47 1.006 ;
        RECT 1.125 0.315 1.215 1.006 ;
        RECT 0.635 0.455 1.215 0.545 ;
        RECT 1.105 0.315 1.215 0.545 ;
        RECT 0.635 0.265 0.725 0.545 ;
        RECT 0.55 0.265 0.725 0.355 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.645 1.096 1.675 1.186 ;
      RECT 1.585 0.863 1.675 1.186 ;
      RECT 1.631 0.838 1.675 1.186 ;
      RECT 0.645 0.675 0.735 1.186 ;
      RECT 1.585 0.863 1.721 0.901 ;
      RECT 1.635 0.23 1.725 0.876 ;
      RECT 0.645 0.675 0.8 0.765 ;
      RECT 1.635 0.23 1.95 0.32 ;
      RECT 0.045 1.04 0.19 1.13 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 0.455 0.445 0.545 0.65 ;
      RECT 0.045 0.445 0.545 0.535 ;
      RECT 0.045 0.23 0.14 0.535 ;
      RECT 0.045 0.23 0.19 0.32 ;
  END
END NOR4BBX1P4H7R

MACRO NOR4BBX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BBX2H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.79 1.08 1.93 1.48 ;
        RECT 0.325 1.07 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.335 -0.08 1.425 0.33 ;
        RECT 0.8 -0.08 0.94 0.305 ;
        RECT 0.325 -0.08 0.415 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.77 0.375 0.95 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.765 0.825 1.945 0.975 ;
      LAYER MET2 ;
        RECT 1.85 0.625 1.95 1.16 ;
      LAYER VIA1 ;
        RECT 1.855 0.855 1.945 0.945 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.845 0.615 0.995 0.795 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.28 0.455 1.575 0.545 ;
        RECT 1.28 0.455 1.37 0.68 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.1 0.855 1.44 0.945 ;
        RECT 1.1 0.395 1.19 0.945 ;
        RECT 0.55 0.395 1.19 0.485 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.665 1.065 1.655 1.155 ;
      RECT 1.565 0.738 1.655 1.155 ;
      RECT 0.665 0.615 0.755 1.155 ;
      RECT 1.611 0.693 1.701 0.776 ;
      RECT 1.655 0.648 1.747 0.73 ;
      RECT 1.655 0.648 1.793 0.684 ;
      RECT 1.701 0.602 1.815 0.65 ;
      RECT 1.747 0.556 1.861 0.616 ;
      RECT 1.793 0.522 1.815 0.65 ;
      RECT 1.815 0.205 1.905 0.571 ;
      RECT 0.045 1.04 0.19 1.13 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 0.045 0.59 0.55 0.68 ;
      RECT 0.045 0.23 0.14 0.68 ;
      RECT 0.045 0.23 0.19 0.32 ;
  END
END NOR4BBX2H7R

MACRO NOR4BBX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BBX3H7R 0 0 ;
  SIZE 3.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.6 1.48 ;
        RECT 1.285 1.21 1.425 1.48 ;
        RECT 0.31 1.205 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.6 0.08 ;
        RECT 3.31 -0.08 3.45 0.305 ;
        RECT 2.81 -0.08 2.95 0.305 ;
        RECT 2.15 -0.08 2.29 0.305 ;
        RECT 1.55 -0.08 1.69 0.305 ;
        RECT 1.045 -0.08 1.135 0.345 ;
        RECT 0.355 -0.08 0.445 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.425 0.57 0.65 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.53 0.35 0.8 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.425 0.62 2.77 0.745 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.93 0.62 3.27 0.745 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.06 0.835 3.545 0.925 ;
        RECT 3.455 0.395 3.545 0.925 ;
        RECT 1.295 0.395 3.545 0.485 ;
        RECT 3.06 0.835 3.2 0.94 ;
        RECT 3.085 0.295 3.175 0.485 ;
        RECT 2.585 0.295 2.675 0.485 ;
        RECT 1.825 0.295 1.915 0.485 ;
        RECT 1.295 0.295 1.385 0.485 ;
      LAYER MET2 ;
        RECT 3.45 0.225 3.55 0.76 ;
      LAYER VIA1 ;
        RECT 3.455 0.455 3.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.31 1.03 3.45 1.12 ;
      RECT 3.31 1.015 3.45 1.12 ;
      RECT 2.81 1.015 2.95 1.12 ;
      RECT 2.31 1.015 2.45 1.12 ;
      RECT 2.56 0.835 2.7 0.94 ;
      RECT 1.8 0.835 1.94 0.94 ;
      RECT 1.8 0.835 2.7 0.925 ;
      RECT 1.045 1.03 2.19 1.12 ;
      RECT 2.05 1.015 2.19 1.12 ;
      RECT 1.55 1.015 1.69 1.12 ;
      RECT 1.045 0.975 1.135 1.12 ;
      RECT 0.07 1.025 0.93 1.115 ;
      RECT 0.84 0.785 0.93 1.115 ;
      RECT 0.07 0.265 0.16 1.115 ;
      RECT 0.84 0.785 1.71 0.875 ;
      RECT 1.62 0.62 1.71 0.875 ;
      RECT 1.62 0.62 2.01 0.71 ;
      RECT 0.575 0.845 0.75 0.935 ;
      RECT 0.66 0.265 0.75 0.935 ;
      RECT 0.66 0.605 1.49 0.695 ;
  END
END NOR4BBX3H7R

MACRO NOR4BBX4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BBX4H7R 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.8 1.48 ;
        RECT 1.335 1.225 1.475 1.48 ;
        RECT 0.315 1.165 0.455 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.8 0.08 ;
        RECT 3.38 -0.08 3.52 0.305 ;
        RECT 2.88 -0.08 3.02 0.305 ;
        RECT 2.2 -0.08 2.34 0.305 ;
        RECT 1.65 -0.08 1.79 0.305 ;
        RECT 1.075 -0.08 1.165 0.345 ;
        RECT 0.355 -0.08 0.445 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.425 0.57 0.66 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.53 0.35 0.8 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.5 0.655 2.84 0.745 ;
      LAYER MET2 ;
        RECT 2.65 0.43 2.75 0.96 ;
      LAYER VIA1 ;
        RECT 2.655 0.655 2.745 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3 0.655 3.34 0.745 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.13 0.885 3.545 0.975 ;
        RECT 3.455 0.395 3.545 0.975 ;
        RECT 1.4 0.395 3.545 0.485 ;
      LAYER MET2 ;
        RECT 3.45 0.625 3.55 1.16 ;
      LAYER VIA1 ;
        RECT 3.455 0.855 3.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.63 0.865 2.77 0.975 ;
      RECT 1.9 0.865 2.77 0.955 ;
      RECT 0.07 0.985 0.93 1.075 ;
      RECT 0.84 0.865 0.93 1.075 ;
      RECT 0.07 0.305 0.16 1.075 ;
      RECT 0.84 0.865 1.77 0.955 ;
      RECT 1.68 0.625 1.77 0.955 ;
      RECT 1.68 0.625 2.11 0.715 ;
      RECT 0.58 0.805 0.75 0.895 ;
      RECT 0.66 0.305 0.75 0.895 ;
      RECT 0.66 0.625 1.54 0.715 ;
      RECT 2.38 1.08 3.52 1.17 ;
      RECT 1.02 1.045 2.29 1.135 ;
  END
END NOR4BBX4H7R

MACRO NOR4BX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BX0P5H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.325 1.025 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.39 -0.08 1.48 0.385 ;
        RECT 0.825 -0.08 0.965 0.175 ;
        RECT 0.31 -0.08 0.45 0.34 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.36 0.825 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.755 0.775 0.98 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.79 0.455 1.06 0.555 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.365 0.625 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.255 1.55 0.785 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.995 1.545 1.175 ;
        RECT 1.15 0.995 1.545 1.085 ;
        RECT 1.15 0.265 1.24 1.085 ;
        RECT 0.56 0.265 1.24 0.355 ;
      LAYER MET2 ;
        RECT 1.45 1.015 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.995 0.19 1.085 ;
      RECT 0.045 0.265 0.135 1.085 ;
      RECT 0.46 0.445 0.55 0.59 ;
      RECT 0.045 0.445 0.55 0.535 ;
      RECT 0.045 0.265 0.14 0.535 ;
      RECT 0.045 0.265 0.19 0.355 ;
  END
END NOR4BX0P5H7R

MACRO NOR4BX0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BX0P7H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.325 1.025 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.39 -0.08 1.48 0.385 ;
        RECT 0.825 -0.08 0.965 0.175 ;
        RECT 0.31 -0.08 0.45 0.34 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.36 0.825 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.728 0.765 0.98 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.455 1.06 0.57 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.365 0.625 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.255 1.55 0.785 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.995 1.545 1.175 ;
        RECT 1.15 0.995 1.545 1.085 ;
        RECT 1.15 0.265 1.24 1.085 ;
        RECT 0.56 0.265 1.24 0.355 ;
      LAYER MET2 ;
        RECT 1.45 1.015 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.995 0.19 1.085 ;
      RECT 0.045 0.265 0.135 1.085 ;
      RECT 0.46 0.445 0.55 0.615 ;
      RECT 0.045 0.445 0.55 0.535 ;
      RECT 0.045 0.265 0.14 0.535 ;
      RECT 0.045 0.265 0.19 0.355 ;
  END
END NOR4BX0P7H7R

MACRO NOR4BX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BX1H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.325 1.025 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.39 -0.08 1.48 0.385 ;
        RECT 0.825 -0.08 0.965 0.175 ;
        RECT 0.31 -0.08 0.45 0.34 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.36 0.825 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.68 0.775 0.98 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.455 1.06 0.6 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.365 0.625 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.255 1.55 0.785 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.995 1.545 1.175 ;
        RECT 1.165 0.995 1.545 1.085 ;
        RECT 1.165 0.265 1.255 1.085 ;
        RECT 0.56 0.265 1.255 0.355 ;
      LAYER MET2 ;
        RECT 1.45 1.015 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.995 0.19 1.085 ;
      RECT 0.045 0.265 0.135 1.085 ;
      RECT 0.455 0.445 0.545 0.65 ;
      RECT 0.045 0.445 0.545 0.535 ;
      RECT 0.045 0.265 0.14 0.535 ;
      RECT 0.045 0.265 0.19 0.355 ;
  END
END NOR4BX1H7R

MACRO NOR4BX1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BX1P4H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.325 1.07 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.39 -0.08 1.48 0.35 ;
        RECT 0.825 -0.08 0.965 0.305 ;
        RECT 0.335 -0.08 0.425 0.345 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.36 0.825 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.64 0.575 0.775 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.855 1.035 0.945 ;
        RECT 0.945 0.706 1.035 0.945 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.365 0.625 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.255 1.55 0.785 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END D
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.995 1.545 1.175 ;
        RECT 1.165 0.995 1.545 1.085 ;
        RECT 1.165 0.34 1.255 1.085 ;
        RECT 0.645 0.395 1.255 0.485 ;
        RECT 1.115 0.34 1.255 0.485 ;
        RECT 0.645 0.265 0.735 0.485 ;
        RECT 0.56 0.265 0.735 0.355 ;
      LAYER MET2 ;
        RECT 1.45 1.015 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Z
  OBS
    LAYER MET1 ;
      RECT 0.045 1.04 0.19 1.13 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 0.455 0.445 0.545 0.65 ;
      RECT 0.045 0.445 0.545 0.535 ;
      RECT 0.045 0.23 0.14 0.535 ;
      RECT 0.045 0.23 0.19 0.32 ;
  END
END NOR4BX1P4H7R

MACRO NOR4BX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BX2H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 0.325 1.07 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.335 -0.08 1.425 0.345 ;
        RECT 0.8 -0.08 0.94 0.305 ;
        RECT 0.325 -0.08 0.415 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.75 0.345 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.62 0.575 0.755 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.855 0.995 0.945 ;
        RECT 0.905 0.615 0.995 0.945 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.28 0.655 1.58 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.1 1.055 1.45 1.145 ;
        RECT 1.1 0.395 1.19 1.145 ;
        RECT 0.575 0.395 1.19 0.485 ;
        RECT 0.575 0.345 0.665 0.485 ;
      LAYER MET2 ;
        RECT 1.25 0.84 1.35 1.22 ;
      LAYER VIA1 ;
        RECT 1.255 1.055 1.345 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 1.06 0.19 1.15 ;
      RECT 0.045 0.23 0.135 1.15 ;
      RECT 0.435 0.565 0.525 0.705 ;
      RECT 0.045 0.565 0.525 0.655 ;
      RECT 0.045 0.23 0.14 0.655 ;
      RECT 0.045 0.23 0.19 0.32 ;
  END
END NOR4BX2H7R

MACRO NOR4BX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BX3H7R 0 0 ;
  SIZE 3 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3 1.48 ;
        RECT 0.8 1.08 0.94 1.48 ;
        RECT 0.325 1.07 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3 0.08 ;
        RECT 2.785 -0.08 2.875 0.345 ;
        RECT 2.285 -0.08 2.375 0.33 ;
        RECT 1.785 -0.08 1.875 0.345 ;
        RECT 1.555 -0.08 1.645 0.345 ;
        RECT 1.055 -0.08 1.145 0.345 ;
        RECT 0.825 -0.08 0.915 0.345 ;
        RECT 0.325 -0.08 0.415 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.62 0.375 0.8 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.15 0.655 1.49 0.745 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.88 0.655 2.22 0.745 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.405 0.655 2.585 0.805 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.51 0.9 2.765 0.99 ;
        RECT 2.675 0.455 2.765 0.99 ;
        RECT 0.645 0.455 2.765 0.545 ;
        RECT 2.51 0.9 2.65 1.02 ;
        RECT 2.535 0.295 2.625 0.545 ;
        RECT 2.035 0.295 2.125 0.545 ;
        RECT 1.305 0.295 1.395 0.545 ;
        RECT 0.645 0.26 0.735 0.545 ;
        RECT 0.55 0.26 0.735 0.35 ;
      LAYER MET2 ;
        RECT 2.25 0.23 2.35 0.76 ;
      LAYER VIA1 ;
        RECT 2.255 0.455 2.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.76 1.11 2.9 1.2 ;
      RECT 2.76 1.08 2.9 1.2 ;
      RECT 2.26 1.095 2.4 1.2 ;
      RECT 1.76 1.08 1.9 1.2 ;
      RECT 2.01 0.885 2.15 1.02 ;
      RECT 1.28 0.885 1.42 1.02 ;
      RECT 1.28 0.885 2.15 0.975 ;
      RECT 1.055 1.11 1.67 1.2 ;
      RECT 1.53 1.08 1.67 1.2 ;
      RECT 1.055 0.9 1.145 1.2 ;
      RECT 0.575 0.9 0.665 1.045 ;
      RECT 0.575 0.9 1.145 0.99 ;
      RECT 0.045 0.96 0.19 1.05 ;
      RECT 0.045 0.29 0.135 1.05 ;
      RECT 0.465 0.64 0.82 0.73 ;
      RECT 0.465 0.44 0.555 0.73 ;
      RECT 0.045 0.44 0.555 0.53 ;
      RECT 0.045 0.29 0.19 0.53 ;
  END
END NOR4BX3H7R

MACRO NOR4BX4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BX4H7R 0 0 ;
  SIZE 3.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.6 1.48 ;
        RECT 0.97 1.08 1.11 1.48 ;
        RECT 0.495 1.07 0.585 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.6 0.08 ;
        RECT 3.185 -0.08 3.275 0.345 ;
        RECT 2.685 -0.08 2.775 0.345 ;
        RECT 2.455 -0.08 2.545 0.345 ;
        RECT 1.955 -0.08 2.045 0.345 ;
        RECT 1.725 -0.08 1.815 0.345 ;
        RECT 1.225 -0.08 1.315 0.345 ;
        RECT 0.995 -0.08 1.085 0.345 ;
        RECT 0.495 -0.08 0.585 0.33 ;
    END
  END VSS
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.395 0.62 0.545 0.8 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.32 0.655 1.66 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.05 0.655 2.39 0.745 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.575 0.655 2.845 0.755 ;
      LAYER MET2 ;
        RECT 2.65 0.43 2.75 0.96 ;
      LAYER VIA1 ;
        RECT 2.655 0.655 2.745 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.935 0.37 3.025 0.95 ;
        RECT 0.815 0.455 3.025 0.545 ;
        RECT 2.205 0.37 2.295 0.545 ;
        RECT 1.475 0.37 1.565 0.545 ;
        RECT 0.815 0.26 0.905 0.545 ;
        RECT 0.72 0.26 0.905 0.35 ;
      LAYER MET2 ;
        RECT 2.85 0.23 2.95 0.76 ;
      LAYER VIA1 ;
        RECT 2.855 0.455 2.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.25 1.065 1.84 1.155 ;
      RECT 1.25 0.9 1.34 1.155 ;
      RECT 0.72 0.9 1.34 0.99 ;
      RECT 0.215 0.92 0.36 1.01 ;
      RECT 0.215 0.33 0.305 1.01 ;
      RECT 0.635 0.64 0.99 0.73 ;
      RECT 0.635 0.44 0.725 0.73 ;
      RECT 0.215 0.44 0.725 0.53 ;
      RECT 0.215 0.33 0.36 0.53 ;
      RECT 2.18 1.08 3.3 1.17 ;
      RECT 1.45 0.885 2.57 0.975 ;
  END
END NOR4BX4H7R

MACRO NOR4X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X0P5H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.07 0.92 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.84 -0.08 0.98 0.175 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.67 0.545 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.65 0.625 0.785 0.825 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.55 1.175 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.6 1.15 1.135 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.875 0.905 1.245 0.995 ;
        RECT 0.045 0.265 1.245 0.355 ;
        RECT 1.025 0.255 1.245 0.355 ;
        RECT 0.875 0.265 0.965 0.995 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.385 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
END NOR4X0P5H7R

MACRO NOR4X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X0P7H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.07 0.952 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.84 -0.08 0.98 0.175 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.67 0.545 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.65 0.595 0.785 0.795 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.55 1.175 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.6 1.15 1.135 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.875 0.905 1.245 0.995 ;
        RECT 0.045 0.265 1.245 0.355 ;
        RECT 1.025 0.255 1.245 0.355 ;
        RECT 0.875 0.265 0.965 0.995 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.385 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
END NOR4X0P7H7R

MACRO NOR4X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X1H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.07 1 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.115 -0.08 1.205 0.2 ;
        RECT 0.585 -0.08 0.675 0.2 ;
        RECT 0.07 -0.08 0.16 0.395 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.62 0.23 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.72 0.545 0.99 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.52 0.78 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.425 1.145 0.725 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.585 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.875 1.055 1.215 1.145 ;
        RECT 0.875 0.315 0.965 1.145 ;
        RECT 0.29 0.315 0.965 0.405 ;
      LAYER MET2 ;
        RECT 1.05 1.015 1.15 1.22 ;
      LAYER VIA1 ;
        RECT 1.055 1.055 1.145 1.145 ;
    END
  END Y
END NOR4X1H7R

MACRO NOR4X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X1P4H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.795 -0.08 0.935 0.305 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.575 0.545 0.8 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.675 0.745 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.575 1.145 0.8 ;
      LAYER MET2 ;
        RECT 1.05 0.6 1.15 1.135 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.845 0.916 1.185 1.006 ;
        RECT 0.07 0.395 1.16 0.485 ;
        RECT 1.055 0.225 1.16 0.485 ;
        RECT 0.845 0.395 0.935 1.006 ;
        RECT 0.57 0.315 0.66 0.485 ;
        RECT 0.07 0.3 0.16 0.485 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.385 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
END NOR4X1P4H7R

MACRO NOR4X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X2H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 0.34 1.055 0.43 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.315 -0.08 1.455 0.305 ;
        RECT 0.815 -0.08 0.955 0.305 ;
        RECT 0.34 -0.08 0.43 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.59 0.545 0.815 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.615 0.76 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.625 1.04 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.195 0.615 1.345 0.795 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.435 0.395 1.545 1.175 ;
        RECT 0.565 0.395 1.545 0.485 ;
      LAYER MET2 ;
        RECT 1.45 0.84 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
END NOR4X2H7R

MACRO NOR4X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X3H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 2.04 -0.08 2.18 0.305 ;
        RECT 1.535 -0.08 1.675 0.305 ;
        RECT 0.795 -0.08 0.935 0.305 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.165 0.655 0.505 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.665 0.655 1.005 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.405 0.655 1.745 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.925 0.655 2.225 0.745 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.04 0.855 2.405 0.945 ;
        RECT 2.315 0.28 2.405 0.945 ;
        RECT 0.07 0.395 2.405 0.485 ;
        RECT 2.04 0.855 2.18 1.02 ;
        RECT 1.81 0.295 1.9 0.485 ;
        RECT 1.07 0.295 1.16 0.485 ;
        RECT 0.57 0.295 0.66 0.485 ;
        RECT 0.07 0.28 0.16 0.485 ;
      LAYER MET2 ;
        RECT 2.25 0.63 2.35 1.16 ;
      LAYER VIA1 ;
        RECT 2.255 0.855 2.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.81 1.11 2.405 1.2 ;
      RECT 2.315 1.055 2.405 1.2 ;
      RECT 1.81 0.915 1.9 1.2 ;
      RECT 1.285 0.915 1.425 1.035 ;
      RECT 1.285 0.915 1.9 1.005 ;
      RECT 0.795 1.125 1.675 1.215 ;
      RECT 1.535 1.095 1.675 1.215 ;
      RECT 0.795 1.095 0.935 1.215 ;
      RECT 0.07 0.915 0.16 1.06 ;
      RECT 0.57 0.915 0.66 1.045 ;
      RECT 1.045 0.915 1.185 1.035 ;
      RECT 0.07 0.915 1.185 1.005 ;
  END
END NOR4X3H7R

MACRO NOR4X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X4H7R 0 0 ;
  SIZE 4.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.2 1.48 ;
        RECT 0.55 1.045 0.69 1.48 ;
        RECT 0.075 1.005 0.165 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.2 0.08 ;
        RECT 3.72 -0.08 3.86 0.175 ;
        RECT 3.19 -0.08 3.33 0.175 ;
        RECT 2.68 -0.08 2.82 0.175 ;
        RECT 2.145 -0.08 2.285 0.175 ;
        RECT 1.63 -0.08 1.77 0.175 ;
        RECT 1.1 -0.08 1.24 0.175 ;
        RECT 0.56 -0.08 0.7 0.175 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.21 0.655 0.75 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.315 0.655 1.855 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.35 0.655 2.89 0.745 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.395 0.635 3.935 0.745 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.475 1.045 4.145 1.135 ;
        RECT 4.025 0.26 4.145 1.135 ;
        RECT 0.295 0.265 4.145 0.355 ;
        RECT 3.985 0.26 4.145 0.355 ;
        RECT 2.945 0.26 3.085 0.355 ;
        RECT 1.895 0.26 2.035 0.355 ;
        RECT 0.825 0.26 0.965 0.355 ;
      LAYER MET2 ;
        RECT 4.05 0.23 4.15 0.76 ;
      LAYER VIA1 ;
        RECT 4.055 0.455 4.145 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.965 0.865 3.055 1.14 ;
      RECT 2.44 0.865 3.865 0.955 ;
      RECT 1.365 1.045 2.83 1.135 ;
      RECT 1.9 0.85 1.99 1.135 ;
      RECT 0.825 0.865 0.915 1.14 ;
      RECT 0.3 0.865 1.755 0.955 ;
  END
END NOR4X4H7R

MACRO NOR4X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X6H7R 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.8 1.48 ;
        RECT 0.84 1.07 0.93 1.48 ;
        RECT 0.34 1.055 0.43 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.8 0.08 ;
        RECT 3.315 -0.08 3.455 0.305 ;
        RECT 2.815 -0.08 2.955 0.305 ;
        RECT 2.315 -0.08 2.455 0.305 ;
        RECT 1.815 -0.08 1.955 0.305 ;
        RECT 1.315 -0.08 1.455 0.305 ;
        RECT 0.815 -0.08 0.955 0.305 ;
        RECT 0.34 -0.08 0.43 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.485 0.655 1.025 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.235 0.655 1.775 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.985 0.655 2.525 0.745 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.71 0.655 3.25 0.745 ;
      LAYER MET2 ;
        RECT 2.85 0.43 2.95 0.96 ;
      LAYER VIA1 ;
        RECT 2.855 0.655 2.945 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.815 1.08 3.575 1.17 ;
        RECT 3.365 1.055 3.575 1.17 ;
        RECT 3.365 0.395 3.455 1.17 ;
        RECT 0.565 0.395 3.455 0.485 ;
      LAYER MET2 ;
        RECT 3.45 0.84 3.55 1.22 ;
      LAYER VIA1 ;
        RECT 3.455 1.055 3.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.065 0.885 3.205 0.975 ;
      RECT 1.315 1.08 2.455 1.17 ;
      RECT 0.565 0.89 1.705 0.98 ;
  END
END NOR4X6H7R

MACRO OA211X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA211X0P5H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.13 1.2 1.28 1.48 ;
        RECT 0.31 1.2 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.29 -0.08 1.38 0.345 ;
        RECT 0.77 -0.08 0.91 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.93 0.455 1.2 0.555 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.675 0.655 0.975 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.445 0.625 0.58 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.625 0.345 0.925 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.54 0.205 1.745 0.375 ;
        RECT 1.48 1.02 1.63 1.16 ;
        RECT 1.54 0.205 1.63 1.16 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.56 ;
      LAYER VIA1 ;
        RECT 1.655 0.255 1.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.23 0.16 1.135 ;
      RECT 0.07 1.02 1.39 1.11 ;
      RECT 1.3 0.73 1.39 1.11 ;
      RECT 0.505 0.265 1.175 0.355 ;
      RECT 1.03 0.255 1.175 0.355 ;
      RECT 0.505 0.26 0.645 0.355 ;
  END
END OA211X0P5H7R

MACRO OA211X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA211X0P7H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.13 1.2 1.28 1.48 ;
        RECT 0.31 1.2 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.29 -0.08 1.38 0.345 ;
        RECT 0.77 -0.08 0.91 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.02 0.455 1.245 0.575 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.675 0.655 0.975 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.445 0.625 0.58 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.625 0.345 0.925 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.54 0.225 1.745 0.375 ;
        RECT 1.48 0.963 1.63 1.103 ;
        RECT 1.54 0.225 1.63 1.103 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.56 ;
      LAYER VIA1 ;
        RECT 1.655 0.255 1.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.23 0.16 1.135 ;
      RECT 0.07 1.02 1.39 1.11 ;
      RECT 1.3 0.73 1.39 1.11 ;
      RECT 0.505 0.265 1.175 0.355 ;
      RECT 1.03 0.255 1.175 0.355 ;
      RECT 0.505 0.255 0.645 0.355 ;
  END
END OA211X0P7H7R

MACRO OA211X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA211X1H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.13 1.2 1.28 1.48 ;
        RECT 0.31 1.2 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.29 -0.08 1.38 0.345 ;
        RECT 0.77 -0.08 0.91 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.02 0.455 1.245 0.575 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.675 0.655 0.975 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.445 0.625 0.58 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.625 0.345 0.925 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.54 0.225 1.745 0.375 ;
        RECT 1.48 0.915 1.63 1.055 ;
        RECT 1.54 0.225 1.63 1.055 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.56 ;
      LAYER VIA1 ;
        RECT 1.655 0.255 1.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.23 0.16 1.135 ;
      RECT 0.07 1.02 1.39 1.11 ;
      RECT 1.3 0.73 1.39 1.11 ;
      RECT 0.505 0.265 1.175 0.355 ;
      RECT 1.03 0.255 1.175 0.355 ;
      RECT 0.505 0.255 0.645 0.355 ;
  END
END OA211X1H7R

MACRO OA211X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA211X1P4H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.13 1.2 1.28 1.48 ;
        RECT 0.31 1.2 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.29 -0.08 1.38 0.345 ;
        RECT 0.77 -0.08 0.91 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.02 0.455 1.245 0.575 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.675 0.655 0.975 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.445 0.625 0.58 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.625 0.345 0.925 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.54 0.225 1.745 0.375 ;
        RECT 1.48 0.891 1.63 1.031 ;
        RECT 1.54 0.225 1.63 1.031 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.56 ;
      LAYER VIA1 ;
        RECT 1.655 0.255 1.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.23 0.16 1.135 ;
      RECT 0.07 1.02 1.345 1.11 ;
      RECT 1.255 0.705 1.345 1.11 ;
      RECT 1.255 0.705 1.45 0.795 ;
      RECT 0.505 0.265 1.175 0.355 ;
      RECT 1.03 0.255 1.175 0.355 ;
      RECT 0.505 0.255 0.645 0.355 ;
  END
END OA211X1P4H7R

MACRO OA211X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA211X2H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.81 1.035 1.9 1.48 ;
        RECT 1.29 1.035 1.38 1.48 ;
        RECT 0.77 1.2 0.91 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.78 -0.08 1.92 0.23 ;
        RECT 1.29 -0.08 1.38 0.435 ;
        RECT 0.31 -0.08 0.45 0.18 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.305 0.455 0.575 0.555 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.655 0.775 0.835 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.93 0.455 1.02 0.65 ;
        RECT 0.825 0.455 1.02 0.545 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.54 0.855 1.945 0.945 ;
        RECT 1.855 0.32 1.945 0.945 ;
        RECT 1.515 0.32 1.945 0.41 ;
        RECT 1.54 0.855 1.63 1.12 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.505 1.02 1.2 1.11 ;
      RECT 1.11 0.25 1.2 1.11 ;
      RECT 1.11 0.675 1.755 0.765 ;
      RECT 1.035 0.25 1.2 0.34 ;
      RECT 0.07 0.275 0.69 0.365 ;
      RECT 0.6 0.225 0.69 0.365 ;
      RECT 0.07 0.225 0.16 0.365 ;
  END
END OA211X2H7R

MACRO OA211X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA211X3H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.81 1.055 1.9 1.48 ;
        RECT 1.29 1.055 1.38 1.48 ;
        RECT 0.77 1.12 0.91 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.79 -0.08 1.88 0.345 ;
        RECT 1.29 -0.08 1.38 0.345 ;
        RECT 0.31 -0.08 0.45 0.18 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.455 0.575 0.545 ;
        RECT 0.425 0.455 0.53 0.675 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.655 0.775 0.835 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.93 0.455 1.02 0.65 ;
        RECT 0.825 0.455 1.02 0.545 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.54 0.855 1.945 0.945 ;
        RECT 1.855 0.495 1.945 0.945 ;
        RECT 1.54 0.495 1.945 0.585 ;
        RECT 1.54 0.855 1.63 1.045 ;
        RECT 1.54 0.295 1.63 0.585 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.505 0.94 1.2 1.03 ;
      RECT 1.11 0.275 1.2 1.03 ;
      RECT 1.11 0.675 1.755 0.765 ;
      RECT 1.035 0.275 1.2 0.365 ;
      RECT 0.045 0.275 0.715 0.365 ;
  END
END OA211X3H7R

MACRO OA211X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA211X4H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.81 1.055 1.9 1.48 ;
        RECT 1.29 1.055 1.38 1.48 ;
        RECT 0.77 1.225 0.91 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.76 -0.08 1.85 0.345 ;
        RECT 1.26 -0.08 1.35 0.345 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.665 0.545 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.64 0.575 0.775 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.855 1.02 0.945 ;
        RECT 0.93 0.665 1.02 0.945 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.515 0.835 1.945 0.925 ;
        RECT 1.855 0.435 1.945 0.925 ;
        RECT 1.51 0.435 1.945 0.525 ;
        RECT 1.51 0.37 1.6 0.525 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.505 1.075 0.649 1.165 ;
      RECT 0.505 1.075 0.651 1.164 ;
      RECT 0.505 1.075 0.689 1.144 ;
      RECT 1.11 0.537 1.2 1.125 ;
      RECT 0.611 1.056 1.2 1.125 ;
      RECT 0.651 1.035 1.2 1.125 ;
      RECT 0.649 1.036 1.2 1.125 ;
      RECT 1.11 0.625 1.755 0.715 ;
      RECT 1.076 0.497 1.166 0.575 ;
      RECT 1.03 0.305 1.12 0.535 ;
      RECT 0.07 0.395 0.66 0.485 ;
      RECT 0.57 0.32 0.66 0.485 ;
      RECT 0.07 0.305 0.16 0.485 ;
  END
END OA211X4H7R

MACRO OA211X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA211X6H7R 0 0 ;
  SIZE 2.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.8 1.48 ;
        RECT 1.795 1.07 1.885 1.48 ;
        RECT 1.295 1.07 1.385 1.48 ;
        RECT 0.585 1.07 0.675 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.8 0.08 ;
        RECT 2 -0.08 2.14 0.305 ;
        RECT 1.525 -0.08 1.615 0.345 ;
        RECT 1.02 -0.08 1.16 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.195 0.595 1.345 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.61 1.005 0.79 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.425 0.755 0.705 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.435 0.565 0.555 0.79 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.275 0.355 2.365 0.945 ;
        RECT 1.635 0.874 2.365 0.945 ;
        RECT 1.674 0.855 2.365 0.945 ;
        RECT 1.75 0.395 2.365 0.485 ;
        RECT 2.045 0.855 2.135 1.17 ;
        RECT 1.545 0.961 1.674 1.003 ;
        RECT 1.591 0.916 1.712 0.964 ;
        RECT 1.545 0.961 1.635 1.13 ;
      LAYER MET2 ;
        RECT 2.05 0.63 2.15 1.16 ;
      LAYER VIA1 ;
        RECT 2.055 0.855 2.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.835 0.88 0.925 1.195 ;
      RECT 0.335 0.88 0.425 1.195 ;
      RECT 0.255 0.88 1.406 0.97 ;
      RECT 0.255 0.88 1.452 0.947 ;
      RECT 1.368 0.861 1.498 0.901 ;
      RECT 0.255 0.38 0.345 0.97 ;
      RECT 1.406 0.819 1.498 0.901 ;
      RECT 1.452 0.773 1.544 0.855 ;
      RECT 1.498 0.727 1.59 0.809 ;
      RECT 1.544 0.681 1.661 0.734 ;
      RECT 1.59 0.641 1.623 0.77 ;
      RECT 1.623 0.625 2.185 0.715 ;
      RECT 0.255 0.38 0.45 0.47 ;
      RECT 0.944 0.395 1.385 0.485 ;
      RECT 1.295 0.345 1.385 0.485 ;
      RECT 0.931 0.35 0.944 0.479 ;
      RECT 0.885 0.321 0.931 0.449 ;
      RECT 0.841 0.19 0.885 0.404 ;
      RECT 0.841 0.376 0.982 0.404 ;
      RECT 0.795 0.19 0.885 0.359 ;
  END
END OA211X6H7R

MACRO OA21X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21X0P5H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.865 1.065 1.155 1.48 ;
        RECT 0.07 0.865 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.045 -0.08 1.185 0.245 ;
        RECT 0.31 -0.08 0.45 0.245 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.575 0.59 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.705 0.655 1.005 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.35 1.025 1.545 1.205 ;
        RECT 1.35 0.31 1.44 1.205 ;
      LAYER MET2 ;
        RECT 1.45 0.84 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.575 0.875 1.205 0.965 ;
      RECT 1.115 0.335 1.205 0.965 ;
      RECT 0.825 0.335 1.205 0.425 ;
      RECT 0.045 0.335 0.715 0.425 ;
  END
END OA21X0P5H7R

MACRO OA21X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21X0P7H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.84 1.055 1.18 1.48 ;
        RECT 0.07 0.865 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.06 -0.08 1.2 0.38 ;
        RECT 0.31 -0.08 0.45 0.245 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.575 0.59 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.705 0.655 0.975 0.755 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.35 1.025 1.545 1.205 ;
        RECT 1.35 0.289 1.44 1.205 ;
      LAYER MET2 ;
        RECT 1.45 0.84 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.575 0.875 1.205 0.965 ;
      RECT 1.115 0.47 1.205 0.965 ;
      RECT 0.955 0.47 1.205 0.56 ;
      RECT 0.94 0.424 0.955 0.553 ;
      RECT 0.896 0.47 1.205 0.523 ;
      RECT 0.85 0.31 0.94 0.478 ;
      RECT 0.85 0.451 0.993 0.478 ;
      RECT 0.045 0.335 0.715 0.425 ;
  END
END OA21X0P7H7R

MACRO OA21X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21X1H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.84 1.055 1.18 1.48 ;
        RECT 0.07 0.865 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.06 -0.08 1.2 0.365 ;
        RECT 0.31 -0.08 0.45 0.245 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.575 0.59 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.705 0.655 1.005 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.35 1.025 1.545 1.205 ;
        RECT 1.35 0.31 1.44 1.205 ;
      LAYER MET2 ;
        RECT 1.45 0.84 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.575 0.875 1.205 0.965 ;
      RECT 1.115 0.475 1.205 0.965 ;
      RECT 0.85 0.475 1.205 0.565 ;
      RECT 0.85 0.31 0.94 0.565 ;
      RECT 0.045 0.335 0.715 0.425 ;
  END
END OA21X1H7R

MACRO OA21X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21X1P4H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.815 1.165 0.955 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.05 -0.08 1.14 0.345 ;
        RECT 0.295 -0.08 0.435 0.325 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.395 0.795 0.545 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.645 0.565 0.765 0.79 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.305 1.415 0.395 ;
        RECT 1.08 0.896 1.345 0.986 ;
        RECT 1.255 0.305 1.345 0.986 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 1.065 0.694 1.155 ;
      RECT 0.55 1.065 0.74 1.132 ;
      RECT 0.656 1.046 0.786 1.086 ;
      RECT 0.694 1.004 0.786 1.086 ;
      RECT 0.74 0.958 0.832 1.04 ;
      RECT 0.786 0.912 0.911 0.961 ;
      RECT 0.832 0.872 0.865 1.001 ;
      RECT 0.865 0.25 0.955 0.916 ;
      RECT 0.865 0.585 1.15 0.675 ;
      RECT 0.795 0.25 0.955 0.34 ;
      RECT 0.07 0.415 0.511 0.505 ;
      RECT 0.07 0.415 0.557 0.482 ;
      RECT 0.473 0.396 0.616 0.423 ;
      RECT 0.557 0.324 0.57 0.453 ;
      RECT 0.07 0.225 0.16 0.505 ;
      RECT 0.511 0.354 0.616 0.423 ;
      RECT 0.57 0.21 0.66 0.378 ;
  END
END OA21X1P4H7R

MACRO OA21X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21X2H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.58 1.185 1.72 1.48 ;
        RECT 1.09 1.035 1.18 1.48 ;
        RECT 0.815 1.185 0.955 1.48 ;
        RECT 0.06 1.075 0.2 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.58 -0.08 1.72 0.215 ;
        RECT 1.09 -0.08 1.18 0.405 ;
        RECT 0.31 -0.08 0.45 0.2 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.045 0.75 0.165 0.975 ;
      LAYER MET2 ;
        RECT 0.05 0.625 0.15 1.16 ;
      LAYER VIA1 ;
        RECT 0.055 0.855 0.145 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.625 0.505 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.65 0.56 0.77 0.785 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.315 1.005 1.745 1.095 ;
        RECT 1.655 0.305 1.745 1.095 ;
        RECT 1.315 0.305 1.745 0.395 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 1.005 0.95 1.095 ;
      RECT 0.86 0.265 0.95 1.095 ;
      RECT 0.86 0.585 1.555 0.675 ;
      RECT 0.045 0.29 0.715 0.38 ;
  END
END OA21X2H7R

MACRO OA21X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21X3H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.325 1.055 1.415 1.48 ;
        RECT 0.825 1.07 0.915 1.48 ;
        RECT 0.06 1.08 0.2 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.55 -0.08 1.64 0.345 ;
        RECT 1.05 -0.08 1.14 0.345 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.695 0.165 0.975 ;
      LAYER MET2 ;
        RECT 0.05 0.625 0.15 1.16 ;
      LAYER VIA1 ;
        RECT 0.055 0.855 0.145 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.625 0.51 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.65 0.555 0.77 0.78 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.115 0.455 1.39 0.545 ;
        RECT 1.3 0.28 1.39 0.545 ;
        RECT 1.05 0.93 1.205 1.02 ;
        RECT 1.115 0.455 1.205 1.02 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.575 0.87 0.665 1.06 ;
      RECT 0.575 0.87 0.95 0.96 ;
      RECT 0.86 0.23 0.95 0.96 ;
      RECT 0.86 0.585 1.025 0.675 ;
      RECT 0.795 0.23 0.95 0.32 ;
      RECT 0.07 0.395 0.576 0.485 ;
      RECT 0.07 0.395 0.622 0.462 ;
      RECT 0.57 0.26 0.66 0.42 ;
      RECT 0.538 0.379 0.66 0.42 ;
      RECT 0.07 0.265 0.16 0.485 ;
  END
END OA21X3H7R

MACRO OA21X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21X4H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.325 1.055 1.415 1.48 ;
        RECT 0.825 1.07 0.915 1.48 ;
        RECT 0.06 1.08 0.2 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.55 -0.08 1.64 0.345 ;
        RECT 1.05 -0.08 1.14 0.345 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.685 0.165 0.975 ;
      LAYER MET2 ;
        RECT 0.05 0.625 0.15 1.16 ;
      LAYER VIA1 ;
        RECT 0.055 0.855 0.145 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.625 0.515 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.65 0.555 0.77 0.78 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.305 1.415 0.395 ;
        RECT 1.05 0.835 1.345 0.925 ;
        RECT 1.255 0.305 1.345 0.925 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.575 0.87 0.665 1.02 ;
      RECT 0.575 0.87 0.95 0.96 ;
      RECT 0.86 0.33 0.95 0.96 ;
      RECT 0.86 0.585 1.055 0.675 ;
      RECT 0.795 0.33 0.95 0.42 ;
      RECT 0.07 0.395 0.581 0.485 ;
      RECT 0.07 0.395 0.627 0.462 ;
      RECT 0.57 0.265 0.66 0.423 ;
      RECT 0.543 0.381 0.66 0.423 ;
      RECT 0.07 0.305 0.16 0.485 ;
  END
END OA21X4H7R

MACRO OA21X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21X6H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 1.545 1.07 1.635 1.48 ;
        RECT 1.045 1.07 1.135 1.48 ;
        RECT 0.265 1.08 0.405 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 1.745 -0.08 1.885 0.305 ;
        RECT 1.27 -0.08 1.36 0.345 ;
        RECT 0.515 -0.08 0.655 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.64 0.365 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.615 0.73 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.85 0.575 0.985 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.495 0.395 2.11 0.485 ;
        RECT 2.02 0.295 2.11 0.485 ;
        RECT 1.795 0.395 1.885 1.165 ;
        RECT 1.295 0.855 1.885 0.945 ;
        RECT 1.295 0.855 1.385 1.195 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.795 0.87 0.885 1.21 ;
      RECT 0.795 0.87 1.165 0.96 ;
      RECT 1.075 0.38 1.165 0.96 ;
      RECT 1.075 0.625 1.675 0.715 ;
      RECT 1.015 0.38 1.165 0.47 ;
      RECT 0.29 0.395 0.905 0.485 ;
      RECT 0.29 0.325 0.38 0.485 ;
  END
END OA21X6H7R

MACRO OA21X8H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21X8H7R 0 0 ;
  SIZE 3.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.4 1.48 ;
        RECT 2.8 1.055 2.89 1.48 ;
        RECT 2.3 1.07 2.39 1.48 ;
        RECT 1.775 1.095 1.915 1.48 ;
        RECT 1.275 1.08 1.415 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.4 0.08 ;
        RECT 2.805 -0.08 2.945 0.305 ;
        RECT 2.305 -0.08 2.445 0.305 ;
        RECT 1.83 -0.08 1.92 0.345 ;
        RECT 0.795 -0.08 0.935 0.305 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.195 0.655 0.535 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.695 0.655 1.035 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.565 0.625 1.745 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.05 0.86 2.945 0.95 ;
        RECT 2.855 0.395 2.945 0.95 ;
        RECT 2.055 0.395 2.945 0.485 ;
        RECT 2.55 0.86 2.64 1.175 ;
        RECT 2.05 0.86 2.14 1.2 ;
      LAYER MET2 ;
        RECT 2.85 0.23 2.95 0.76 ;
      LAYER VIA1 ;
        RECT 2.855 0.455 2.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.525 0.9 1.665 0.995 ;
      RECT 0.795 0.9 0.935 0.995 ;
      RECT 0.795 0.9 1.788 0.99 ;
      RECT 0.795 0.9 1.834 0.967 ;
      RECT 1.75 0.881 1.88 0.921 ;
      RECT 1.31 0.36 1.4 0.99 ;
      RECT 1.788 0.839 1.88 0.921 ;
      RECT 1.834 0.793 1.926 0.875 ;
      RECT 1.88 0.747 1.972 0.829 ;
      RECT 1.88 0.747 2.018 0.783 ;
      RECT 1.926 0.701 2.025 0.757 ;
      RECT 1.926 0.701 2.063 0.734 ;
      RECT 2.025 0.625 2.765 0.715 ;
      RECT 1.972 0.655 2.765 0.715 ;
      RECT 2.018 0.628 2.025 0.757 ;
      RECT 1.31 0.36 1.45 0.45 ;
      RECT 0.07 0.395 1.16 0.485 ;
      RECT 1.07 0.17 1.16 0.485 ;
      RECT 0.57 0.32 0.66 0.485 ;
      RECT 0.07 0.305 0.16 0.485 ;
      RECT 1.6 0.17 1.69 0.345 ;
      RECT 1.07 0.17 1.69 0.26 ;
      RECT 0.57 1.085 1.185 1.175 ;
      RECT 1.045 1.08 1.185 1.175 ;
      RECT 0.57 0.905 0.66 1.175 ;
      RECT 0.07 0.905 0.16 1.045 ;
      RECT 0.07 0.905 0.66 0.995 ;
  END
END OA21X8H7R

MACRO OA221X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA221X0P5H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.58 1.07 1.67 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.58 -0.08 1.67 0.33 ;
        RECT 1.055 -0.08 1.195 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.015 0.845 1.285 0.945 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.395 0.595 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.71 0.645 0.98 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.59 0.585 0.79 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.425 0.345 0.65 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.805 1.04 1.945 1.13 ;
        RECT 1.855 0.23 1.945 1.13 ;
        RECT 1.805 0.23 1.945 0.32 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.525 1.055 1.465 1.145 ;
      RECT 1.375 0.865 1.465 1.145 ;
      RECT 0.045 0.915 0.185 1.13 ;
      RECT 0.525 0.915 0.615 1.145 ;
      RECT 0.045 0.915 0.615 1.005 ;
      RECT 1.375 0.865 1.765 0.955 ;
      RECT 1.675 0.805 1.765 0.955 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.56 0.41 1.42 0.5 ;
      RECT 1.33 0.22 1.42 0.5 ;
      RECT 0.56 0.35 0.7 0.5 ;
      RECT 0.32 0.17 0.41 0.33 ;
      RECT 0.825 0.17 0.965 0.32 ;
      RECT 0.32 0.17 0.965 0.26 ;
  END
END OA221X0P5H7R

MACRO OA221X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA221X0P7H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.58 1.07 1.67 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.58 -0.08 1.67 0.33 ;
        RECT 1.055 -0.08 1.195 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1 0.845 1.27 0.945 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.395 0.595 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.715 0.645 0.985 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.59 0.59 0.79 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.42 0.345 0.645 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.805 1.04 1.945 1.13 ;
        RECT 1.855 0.23 1.945 1.13 ;
        RECT 1.805 0.23 1.945 0.32 ;
      LAYER MET2 ;
        RECT 1.85 0.225 1.95 0.76 ;
      LAYER VIA1 ;
        RECT 1.855 0.455 1.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.525 1.055 1.465 1.145 ;
      RECT 1.375 0.865 1.465 1.145 ;
      RECT 0.045 0.915 0.185 1.13 ;
      RECT 0.525 0.915 0.615 1.145 ;
      RECT 0.045 0.915 0.615 1.005 ;
      RECT 1.375 0.865 1.765 0.955 ;
      RECT 1.675 0.77 1.765 0.955 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.56 0.41 1.42 0.5 ;
      RECT 1.33 0.22 1.42 0.5 ;
      RECT 0.56 0.35 0.7 0.5 ;
      RECT 0.32 0.17 0.41 0.33 ;
      RECT 0.825 0.17 0.965 0.32 ;
      RECT 0.32 0.17 0.965 0.26 ;
  END
END OA221X0P7H7R

MACRO OA221X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA221X1H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.58 1.07 1.67 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.58 -0.08 1.67 0.33 ;
        RECT 1.055 -0.08 1.195 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.005 0.845 1.275 0.945 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.395 0.595 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.71 0.645 0.98 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.59 0.585 0.79 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.425 0.345 0.65 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.805 0.96 1.945 1.05 ;
        RECT 1.855 0.23 1.945 1.05 ;
        RECT 1.805 0.23 1.945 0.32 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.525 1.055 1.465 1.145 ;
      RECT 1.375 0.865 1.465 1.145 ;
      RECT 0.045 0.915 0.185 1.13 ;
      RECT 0.525 0.915 0.615 1.145 ;
      RECT 0.045 0.915 0.615 1.005 ;
      RECT 1.375 0.865 1.679 0.955 ;
      RECT 1.375 0.865 1.725 0.932 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 1.675 0.725 1.765 0.889 ;
      RECT 1.641 0.848 1.765 0.889 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.56 0.41 1.42 0.5 ;
      RECT 1.33 0.22 1.42 0.5 ;
      RECT 0.56 0.35 0.7 0.5 ;
      RECT 0.32 0.17 0.41 0.33 ;
      RECT 0.825 0.17 0.965 0.32 ;
      RECT 0.32 0.17 0.965 0.26 ;
  END
END OA221X1H7R

MACRO OA221X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA221X1P4H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.58 1.07 1.67 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.58 -0.08 1.67 0.33 ;
        RECT 1.055 -0.08 1.195 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.995 0.845 1.265 0.945 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.395 0.595 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.705 0.645 0.975 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.59 0.585 0.79 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.425 0.345 0.65 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.805 0.916 1.945 1.006 ;
        RECT 1.855 0.326 1.945 1.006 ;
        RECT 1.805 0.326 1.945 0.416 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.525 1.055 1.465 1.145 ;
      RECT 1.375 0.865 1.465 1.145 ;
      RECT 0.045 0.915 0.185 1.13 ;
      RECT 0.525 0.915 0.615 1.145 ;
      RECT 0.045 0.915 0.615 1.005 ;
      RECT 1.375 0.865 1.632 0.955 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 1.675 0.681 1.721 0.889 ;
      RECT 1.594 0.846 1.721 0.889 ;
      RECT 1.632 0.805 1.675 0.934 ;
      RECT 1.675 0.681 1.765 0.844 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.56 0.41 1.42 0.5 ;
      RECT 1.33 0.22 1.42 0.5 ;
      RECT 0.56 0.35 0.7 0.5 ;
      RECT 0.32 0.17 0.41 0.33 ;
      RECT 0.825 0.17 0.965 0.32 ;
      RECT 0.32 0.17 0.965 0.26 ;
  END
END OA221X1P4H7R

MACRO OA221X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA221X2H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 1.58 1.07 1.67 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 1.58 -0.08 1.67 0.33 ;
        RECT 1.055 -0.08 1.195 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.995 0.845 1.265 0.945 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.395 0.595 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.705 0.645 0.975 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.59 0.585 0.79 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.425 0.345 0.65 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.805 0.905 1.945 0.995 ;
        RECT 1.855 0.38 1.945 0.995 ;
        RECT 1.805 0.38 1.945 0.47 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.525 1.065 1.465 1.155 ;
      RECT 1.375 0.865 1.465 1.155 ;
      RECT 0.045 0.915 0.185 1.13 ;
      RECT 0.525 0.915 0.615 1.155 ;
      RECT 0.045 0.915 0.615 1.005 ;
      RECT 1.375 0.865 1.624 0.955 ;
      RECT 1.375 0.865 1.67 0.932 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 1.586 0.846 1.721 0.881 ;
      RECT 1.67 0.778 1.675 0.907 ;
      RECT 1.624 0.804 1.721 0.881 ;
      RECT 1.675 0.615 1.765 0.836 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.56 0.41 1.42 0.5 ;
      RECT 1.33 0.22 1.42 0.5 ;
      RECT 0.56 0.35 0.7 0.5 ;
      RECT 0.32 0.17 0.41 0.33 ;
      RECT 0.825 0.17 0.965 0.32 ;
      RECT 0.32 0.17 0.965 0.26 ;
  END
END OA221X2H7R

MACRO OA221X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA221X3H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 2.08 1.055 2.17 1.48 ;
        RECT 1.58 1.07 1.67 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 2.08 -0.08 2.17 0.345 ;
        RECT 1.58 -0.08 1.67 0.33 ;
        RECT 1.055 -0.08 1.195 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.855 1.24 0.945 ;
        RECT 1.15 0.745 1.24 0.945 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.395 0.595 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.715 0.645 0.985 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.59 0.585 0.79 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.425 0.345 0.65 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.805 0.94 1.945 1.03 ;
        RECT 1.855 0.32 1.945 1.03 ;
        RECT 1.805 0.32 1.945 0.41 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.525 1.035 1.465 1.125 ;
      RECT 1.375 0.865 1.465 1.125 ;
      RECT 0.045 0.915 0.185 1.05 ;
      RECT 0.525 0.915 0.615 1.125 ;
      RECT 0.045 0.915 0.615 1.005 ;
      RECT 1.375 0.865 1.662 0.955 ;
      RECT 1.375 0.865 1.721 0.919 ;
      RECT 0.045 0.25 0.135 1.05 ;
      RECT 1.675 0.71 1.765 0.874 ;
      RECT 1.624 0.846 1.765 0.874 ;
      RECT 1.662 0.82 1.675 0.949 ;
      RECT 0.045 0.25 0.185 0.34 ;
      RECT 0.56 0.41 1.42 0.5 ;
      RECT 1.33 0.28 1.42 0.5 ;
      RECT 0.56 0.35 0.7 0.5 ;
      RECT 0.32 0.17 0.41 0.33 ;
      RECT 0.825 0.17 0.965 0.32 ;
      RECT 0.32 0.17 0.965 0.26 ;
  END
END OA221X3H7R

MACRO OA221X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA221X4H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 2.08 0.855 2.17 1.48 ;
        RECT 1.58 1.07 1.67 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 2.08 -0.08 2.17 0.345 ;
        RECT 1.58 -0.08 1.67 0.33 ;
        RECT 1.055 -0.08 1.195 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.855 1.24 0.945 ;
        RECT 1.15 0.71 1.24 0.945 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.395 0.595 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.705 0.645 0.975 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.59 0.585 0.79 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.425 0.345 0.655 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.805 0.9 1.945 0.99 ;
        RECT 1.855 0.395 1.945 0.99 ;
        RECT 1.805 0.395 1.945 0.485 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.525 1.035 1.465 1.125 ;
      RECT 1.375 0.865 1.465 1.125 ;
      RECT 0.525 0.915 0.615 1.125 ;
      RECT 0.045 0.915 0.185 1.01 ;
      RECT 0.045 0.915 0.615 1.005 ;
      RECT 1.375 0.865 1.622 0.955 ;
      RECT 1.375 0.865 1.668 0.932 ;
      RECT 0.045 0.25 0.135 1.01 ;
      RECT 1.584 0.846 1.721 0.879 ;
      RECT 1.668 0.777 1.675 0.906 ;
      RECT 1.622 0.804 1.721 0.879 ;
      RECT 1.675 0.615 1.765 0.834 ;
      RECT 0.045 0.25 0.185 0.34 ;
      RECT 0.56 0.41 1.42 0.5 ;
      RECT 1.33 0.32 1.42 0.5 ;
      RECT 0.56 0.36 0.7 0.5 ;
      RECT 0.32 0.17 0.41 0.33 ;
      RECT 0.825 0.17 0.965 0.32 ;
      RECT 0.32 0.17 0.965 0.26 ;
  END
END OA221X4H7R

MACRO OA222X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA222X0P5H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 1.86 1.07 1.95 1.48 ;
        RECT 1.105 1.225 1.245 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 1.86 -0.08 1.95 0.33 ;
        RECT 1.335 -0.08 1.475 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.65 0.595 1.8 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.35 0.83 1.575 0.95 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.95 0.835 1.175 0.955 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.71 0.645 0.98 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.505 0.855 0.775 0.945 ;
        RECT 0.505 0.805 0.595 0.945 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.085 1.04 2.235 1.13 ;
        RECT 2.145 0.225 2.235 1.13 ;
        RECT 2.055 0.225 2.235 0.375 ;
      LAYER MET2 ;
        RECT 2.05 0.18 2.15 0.56 ;
      LAYER VIA1 ;
        RECT 2.055 0.255 2.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.325 1.045 1.77 1.135 ;
      RECT 1.68 0.865 1.77 1.135 ;
      RECT 0.325 0.35 0.415 1.135 ;
      RECT 1.68 0.865 2.05 0.955 ;
      RECT 1.96 0.805 2.05 0.955 ;
      RECT 0.31 0.35 0.45 0.44 ;
      RECT 0.84 0.41 1.7 0.5 ;
      RECT 1.61 0.22 1.7 0.5 ;
      RECT 0.84 0.35 0.98 0.5 ;
      RECT 0.07 0.17 0.16 0.345 ;
      RECT 0.6 0.17 0.69 0.33 ;
      RECT 1.105 0.17 1.245 0.32 ;
      RECT 0.07 0.17 1.245 0.26 ;
  END
END OA222X0P5H7R

MACRO OA222X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA222X0P7H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 1.86 1.07 1.95 1.48 ;
        RECT 1.105 1.225 1.245 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 1.86 -0.08 1.95 0.33 ;
        RECT 1.335 -0.08 1.475 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.625 0.595 1.805 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.35 0.83 1.575 0.95 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.96 0.835 1.185 0.955 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.705 0.645 0.975 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.505 0.855 0.775 0.945 ;
        RECT 0.505 0.805 0.595 0.945 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.085 1.01 2.235 1.1 ;
        RECT 2.145 0.225 2.235 1.1 ;
        RECT 2.055 0.225 2.235 0.375 ;
      LAYER MET2 ;
        RECT 2.05 0.18 2.15 0.56 ;
      LAYER VIA1 ;
        RECT 2.055 0.255 2.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.325 1.045 1.755 1.135 ;
      RECT 1.665 0.835 1.755 1.135 ;
      RECT 0.325 0.35 0.415 1.135 ;
      RECT 1.665 0.835 2.055 0.925 ;
      RECT 1.965 0.77 2.055 0.925 ;
      RECT 0.31 0.35 0.45 0.44 ;
      RECT 0.84 0.41 1.7 0.5 ;
      RECT 1.61 0.22 1.7 0.5 ;
      RECT 0.84 0.35 0.98 0.5 ;
      RECT 0.07 0.17 0.16 0.345 ;
      RECT 0.6 0.17 0.69 0.33 ;
      RECT 1.105 0.17 1.245 0.32 ;
      RECT 0.07 0.17 1.245 0.26 ;
  END
END OA222X0P7H7R

MACRO OA222X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA222X1H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 1.92 1.215 2.06 1.48 ;
        RECT 1.095 1.215 1.235 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 1.935 -0.08 2.075 0.34 ;
        RECT 0.295 -0.08 0.435 0.325 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.42 0.855 0.59 0.945 ;
        RECT 0.42 0.725 0.51 0.945 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.825 1.05 0.945 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.6 0.595 0.78 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.225 0.825 1.45 0.945 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.595 0.625 1.745 0.805 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.24 0.25 2.345 1.13 ;
      LAYER MET2 ;
        RECT 2.25 0.23 2.35 0.76 ;
      LAYER VIA1 ;
        RECT 2.255 0.455 2.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.545 1.035 1.925 1.125 ;
      RECT 1.835 0.445 1.925 1.125 ;
      RECT 1.835 0.57 2.145 0.66 ;
      RECT 1.385 0.445 1.475 0.645 ;
      RECT 1.385 0.445 1.925 0.535 ;
      RECT 1.66 0.205 1.75 0.535 ;
      RECT 1.135 0.23 1.225 0.63 ;
      RECT 0.795 0.23 1.225 0.325 ;
      RECT 0.795 0.23 1.525 0.32 ;
      RECT 0.885 0.415 0.975 0.63 ;
      RECT 0.07 0.415 0.975 0.505 ;
      RECT 0.57 0.24 0.66 0.505 ;
      RECT 0.07 0.225 0.16 0.505 ;
  END
END OA222X1H7R

MACRO OA222X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA222X1P4H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 1.86 1.07 1.95 1.48 ;
        RECT 1.105 1.225 1.245 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 1.86 -0.08 1.95 0.33 ;
        RECT 1.335 -0.08 1.475 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.62 0.595 1.8 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.35 0.83 1.575 0.95 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.955 0.835 1.18 0.955 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.71 0.645 0.98 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.505 0.855 0.775 0.945 ;
        RECT 0.505 0.805 0.595 0.945 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.085 1.01 2.235 1.1 ;
        RECT 2.145 0.225 2.235 1.1 ;
        RECT 2.055 0.225 2.235 0.375 ;
      LAYER MET2 ;
        RECT 2.05 0.18 2.15 0.56 ;
      LAYER VIA1 ;
        RECT 2.055 0.255 2.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.325 1.045 1.77 1.135 ;
      RECT 1.68 0.835 1.77 1.135 ;
      RECT 0.325 0.35 0.415 1.135 ;
      RECT 1.68 0.835 2.055 0.925 ;
      RECT 1.965 0.68 2.055 0.925 ;
      RECT 0.31 0.35 0.45 0.44 ;
      RECT 0.84 0.41 1.7 0.5 ;
      RECT 1.61 0.22 1.7 0.5 ;
      RECT 0.84 0.35 0.98 0.5 ;
      RECT 0.07 0.17 0.16 0.345 ;
      RECT 0.6 0.17 0.69 0.33 ;
      RECT 1.105 0.17 1.245 0.32 ;
      RECT 0.07 0.17 1.245 0.26 ;
  END
END OA222X1P4H7R

MACRO OA222X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA222X2H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 1.92 1.07 2.01 1.48 ;
        RECT 1.105 1.225 1.245 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 1.92 -0.08 2.01 0.33 ;
        RECT 1.395 -0.08 1.535 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.77 0.595 1.975 0.745 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.41 0.83 1.635 0.95 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.955 0.835 1.18 0.955 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.685 0.645 0.975 0.745 ;
        RECT 0.685 0.645 0.865 0.765 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.505 0.855 0.775 0.945 ;
        RECT 0.505 0.805 0.595 0.945 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.115 1.025 2.375 1.175 ;
        RECT 2.25 0.38 2.375 1.175 ;
        RECT 2.145 0.38 2.375 0.47 ;
      LAYER MET2 ;
        RECT 2.25 0.84 2.35 1.22 ;
      LAYER VIA1 ;
        RECT 2.255 1.055 2.345 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.325 1.045 1.815 1.135 ;
      RECT 1.725 0.835 1.815 1.135 ;
      RECT 0.325 0.35 0.415 1.135 ;
      RECT 1.725 0.835 2.16 0.925 ;
      RECT 2.07 0.615 2.16 0.925 ;
      RECT 0.31 0.35 0.45 0.44 ;
      RECT 1.111 0.54 1.429 0.63 ;
      RECT 1.082 0.487 1.111 0.616 ;
      RECT 1.036 0.45 1.082 0.578 ;
      RECT 1.391 0.521 1.506 0.576 ;
      RECT 1.429 0.486 1.46 0.615 ;
      RECT 1.036 0.521 1.149 0.578 ;
      RECT 0.99 0.404 1.036 0.532 ;
      RECT 1.46 0.41 1.552 0.53 ;
      RECT 0.981 0.487 1.111 0.505 ;
      RECT 1.429 0.486 1.559 0.504 ;
      RECT 1.67 0.22 1.76 0.5 ;
      RECT 0.84 0.35 0.99 0.5 ;
      RECT 1.46 0.41 1.76 0.5 ;
      RECT 1.19 0.17 1.28 0.45 ;
      RECT 0.6 0.17 0.69 0.45 ;
      RECT 0.07 0.17 0.16 0.45 ;
      RECT 0.07 0.17 1.28 0.26 ;
  END
END OA222X2H7R

MACRO OA222X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA222X3H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 2.375 1.055 2.465 1.48 ;
        RECT 1.875 1.07 1.965 1.48 ;
        RECT 1.105 1.225 1.245 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 2.375 -0.08 2.465 0.345 ;
        RECT 1.875 -0.08 1.965 0.33 ;
        RECT 1.35 -0.08 1.49 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.655 0.625 1.89 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.425 0.855 1.59 0.945 ;
        RECT 1.425 0.725 1.555 0.945 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.855 1.18 0.95 ;
        RECT 1.035 0.77 1.18 0.95 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.625 0.945 0.775 ;
        RECT 0.74 0.625 0.945 0.765 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.505 0.855 0.775 0.945 ;
        RECT 0.505 0.725 0.595 0.945 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.055 1.025 2.25 1.175 ;
        RECT 2.16 0.32 2.25 1.175 ;
        RECT 2.1 0.32 2.25 0.41 ;
      LAYER MET2 ;
        RECT 2.05 0.84 2.15 1.22 ;
      LAYER VIA1 ;
        RECT 2.055 1.055 2.145 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.325 1.045 1.77 1.135 ;
      RECT 1.68 0.865 1.77 1.135 ;
      RECT 0.325 0.35 0.415 1.135 ;
      RECT 1.68 0.865 1.989 0.955 ;
      RECT 1.68 0.865 2.035 0.932 ;
      RECT 1.98 0.71 2.07 0.892 ;
      RECT 1.951 0.85 2.07 0.892 ;
      RECT 0.31 0.35 0.45 0.44 ;
      RECT 0.84 0.44 1.715 0.53 ;
      RECT 1.625 0.28 1.715 0.53 ;
      RECT 0.84 0.35 0.98 0.53 ;
      RECT 0.07 0.17 0.16 0.39 ;
      RECT 0.6 0.17 0.69 0.375 ;
      RECT 1.105 0.17 1.245 0.35 ;
      RECT 0.07 0.17 1.245 0.26 ;
  END
END OA222X3H7R

MACRO OA222X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA222X4H7R 0 0 ;
  SIZE 2.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.8 1.48 ;
        RECT 2.335 1.08 2.475 1.48 ;
        RECT 1.86 1.07 1.95 1.48 ;
        RECT 1.105 1.225 1.245 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.8 0.08 ;
        RECT 2.36 -0.08 2.45 0.345 ;
        RECT 1.86 -0.08 1.95 0.33 ;
        RECT 1.335 -0.08 1.475 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.655 0.595 1.805 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.42 0.855 1.575 0.945 ;
        RECT 1.42 0.735 1.56 0.945 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.855 1.175 0.945 ;
        RECT 1.035 0.735 1.175 0.945 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.625 0.945 0.775 ;
        RECT 0.735 0.625 0.945 0.765 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.505 0.855 0.775 0.945 ;
        RECT 0.505 0.685 0.595 0.945 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.085 0.885 2.345 0.975 ;
        RECT 2.145 0.825 2.345 0.975 ;
        RECT 2.145 0.395 2.235 0.975 ;
        RECT 2.085 0.395 2.235 0.485 ;
      LAYER MET2 ;
        RECT 2.25 0.63 2.35 1.16 ;
      LAYER VIA1 ;
        RECT 2.255 0.855 2.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.325 1.045 1.755 1.135 ;
      RECT 1.665 0.865 1.755 1.135 ;
      RECT 0.325 0.35 0.415 1.135 ;
      RECT 1.665 0.865 1.882 0.955 ;
      RECT 1.665 0.865 1.928 0.932 ;
      RECT 1.844 0.846 1.965 0.891 ;
      RECT 1.882 0.804 2.011 0.849 ;
      RECT 1.928 0.762 1.965 0.891 ;
      RECT 1.965 0.615 2.055 0.804 ;
      RECT 0.31 0.35 0.45 0.44 ;
      RECT 0.84 0.415 1.7 0.505 ;
      RECT 1.61 0.22 1.7 0.505 ;
      RECT 0.84 0.35 0.98 0.505 ;
      RECT 0.07 0.17 0.16 0.35 ;
      RECT 0.6 0.17 0.69 0.335 ;
      RECT 1.105 0.17 1.245 0.325 ;
      RECT 0.07 0.17 1.245 0.26 ;
  END
END OA222X4H7R

MACRO OA22X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22X0P5H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.07 1.07 1.16 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.36 -0.08 1.45 0.345 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.595 0.545 0.795 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.565 1.175 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.635 0.75 0.755 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.335 1.055 1.7 1.145 ;
        RECT 1.61 0.205 1.7 1.145 ;
      LAYER MET2 ;
        RECT 1.45 0.84 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.545 1.065 0.935 1.155 ;
      RECT 0.845 0.35 0.935 1.155 ;
      RECT 0.845 0.85 1.38 0.94 ;
      RECT 1.29 0.8 1.38 0.94 ;
      RECT 0.825 0.35 0.965 0.44 ;
      RECT 0.07 0.395 0.66 0.485 ;
      RECT 0.57 0.17 0.66 0.485 ;
      RECT 0.07 0.205 0.16 0.485 ;
      RECT 1.13 0.17 1.22 0.345 ;
      RECT 0.57 0.17 1.22 0.26 ;
  END
END OA22X0P5H7R

MACRO OA22X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22X0P7H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.07 1.07 1.16 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.36 -0.08 1.45 0.345 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.595 0.545 0.795 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.565 1.175 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.635 0.75 0.755 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.335 1.055 1.7 1.145 ;
        RECT 1.61 0.205 1.7 1.145 ;
      LAYER MET2 ;
        RECT 1.45 0.84 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.545 1.065 0.935 1.155 ;
      RECT 0.845 0.35 0.935 1.155 ;
      RECT 0.845 0.835 1.38 0.925 ;
      RECT 1.29 0.785 1.38 0.925 ;
      RECT 0.825 0.35 0.965 0.44 ;
      RECT 0.07 0.395 0.66 0.485 ;
      RECT 0.57 0.17 0.66 0.485 ;
      RECT 0.07 0.205 0.16 0.485 ;
      RECT 1.13 0.17 1.22 0.345 ;
      RECT 0.57 0.17 1.22 0.26 ;
  END
END OA22X0P7H7R

MACRO OA22X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22X1H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.07 1.07 1.16 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.36 -0.08 1.45 0.345 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.595 0.545 0.795 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.565 1.175 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.635 0.75 0.755 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.335 1.055 1.7 1.145 ;
        RECT 1.61 0.265 1.7 1.145 ;
      LAYER MET2 ;
        RECT 1.45 0.84 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.545 1.065 0.935 1.155 ;
      RECT 0.845 0.35 0.935 1.155 ;
      RECT 0.845 0.835 1.38 0.925 ;
      RECT 1.29 0.75 1.38 0.925 ;
      RECT 0.825 0.35 0.965 0.44 ;
      RECT 0.07 0.395 0.66 0.485 ;
      RECT 0.57 0.17 0.66 0.485 ;
      RECT 0.07 0.205 0.16 0.485 ;
      RECT 1.13 0.17 1.22 0.345 ;
      RECT 0.57 0.17 1.22 0.26 ;
  END
END OA22X1H7R

MACRO OA22X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22X1P4H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.07 1.07 1.16 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.36 -0.08 1.45 0.345 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.595 0.545 0.795 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.565 1.175 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.635 0.75 0.755 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.335 1.055 1.7 1.145 ;
        RECT 1.61 0.301 1.7 1.145 ;
      LAYER MET2 ;
        RECT 1.45 0.84 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.545 1.065 0.935 1.155 ;
      RECT 0.845 0.35 0.935 1.155 ;
      RECT 0.845 0.845 1.38 0.935 ;
      RECT 1.29 0.705 1.38 0.935 ;
      RECT 0.825 0.35 0.965 0.44 ;
      RECT 0.07 0.395 0.66 0.485 ;
      RECT 0.57 0.17 0.66 0.485 ;
      RECT 0.07 0.205 0.16 0.485 ;
      RECT 1.13 0.17 1.22 0.345 ;
      RECT 0.57 0.17 1.22 0.26 ;
  END
END OA22X1P4H7R

MACRO OA22X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22X2H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.07 1.07 1.16 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.36 -0.08 1.45 0.345 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.595 0.545 0.795 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.03 0.55 1.15 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.64 0.75 0.76 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.335 1.055 1.7 1.145 ;
        RECT 1.61 0.29 1.7 1.145 ;
      LAYER MET2 ;
        RECT 1.45 0.84 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.545 1.065 0.94 1.155 ;
      RECT 0.85 0.35 0.94 1.155 ;
      RECT 0.85 0.865 1.38 0.955 ;
      RECT 1.29 0.64 1.38 0.955 ;
      RECT 0.825 0.35 0.965 0.44 ;
      RECT 0.07 0.395 0.66 0.485 ;
      RECT 0.57 0.17 0.66 0.485 ;
      RECT 0.07 0.205 0.16 0.485 ;
      RECT 1.13 0.17 1.22 0.345 ;
      RECT 0.57 0.17 1.22 0.26 ;
  END
END OA22X2H7R

MACRO OA22X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22X3H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.65 1.225 1.79 1.48 ;
        RECT 1.07 1.07 1.16 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.86 -0.08 1.95 0.345 ;
        RECT 1.36 -0.08 1.45 0.345 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.595 0.545 0.795 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.565 1.175 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.705 0.755 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.61 0.295 1.7 1.046 ;
        RECT 1.541 1.036 1.656 1.091 ;
        RECT 1.579 1.001 1.61 1.13 ;
        RECT 1.335 1.055 1.579 1.145 ;
      LAYER MET2 ;
        RECT 1.45 0.84 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.545 1.065 0.935 1.155 ;
      RECT 0.845 0.35 0.935 1.155 ;
      RECT 0.845 0.835 1.38 0.925 ;
      RECT 1.29 0.735 1.38 0.925 ;
      RECT 0.825 0.35 0.965 0.44 ;
      RECT 0.07 0.395 0.66 0.485 ;
      RECT 0.57 0.17 0.66 0.485 ;
      RECT 0.07 0.205 0.16 0.485 ;
      RECT 1.13 0.17 1.22 0.345 ;
      RECT 0.57 0.17 1.22 0.26 ;
  END
END OA22X3H7R

MACRO OA22X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22X4H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 1.65 1.205 1.79 1.48 ;
        RECT 1.07 1.07 1.16 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 1.86 -0.08 1.95 0.345 ;
        RECT 1.36 -0.08 1.45 0.345 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.595 0.545 0.795 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.015 0.595 1.195 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.675 0.745 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.61 0.37 1.7 1.046 ;
        RECT 1.541 1.036 1.656 1.091 ;
        RECT 1.579 1.001 1.61 1.13 ;
        RECT 1.335 1.055 1.579 1.145 ;
      LAYER MET2 ;
        RECT 1.45 0.84 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.545 1.065 0.925 1.155 ;
      RECT 0.835 0.35 0.925 1.155 ;
      RECT 0.835 0.835 1.38 0.925 ;
      RECT 1.29 0.64 1.38 0.925 ;
      RECT 0.825 0.35 0.965 0.44 ;
      RECT 0.07 0.395 0.66 0.485 ;
      RECT 0.57 0.17 0.66 0.485 ;
      RECT 0.07 0.305 0.16 0.485 ;
      RECT 1.13 0.17 1.22 0.345 ;
      RECT 0.57 0.17 1.22 0.26 ;
  END
END OA22X4H7R

MACRO OA22X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22X6H7R 0 0 ;
  SIZE 2.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.8 1.48 ;
        RECT 1.902 1.225 2.042 1.48 ;
        RECT 1.322 1.07 1.412 1.48 ;
        RECT 0.322 1.055 0.412 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.8 0.08 ;
        RECT 2.027 -0.08 2.167 0.305 ;
        RECT 1.552 -0.08 1.642 0.345 ;
        RECT 0.547 -0.08 0.687 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.595 0.545 0.795 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.615 0.745 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.282 0.605 1.575 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.615 1.005 0.795 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.777 0.395 2.392 0.485 ;
        RECT 2.302 0.345 2.392 0.485 ;
        RECT 2.242 0.395 2.345 1.175 ;
        RECT 1.587 1.02 2.345 1.11 ;
      LAYER MET2 ;
        RECT 2.25 0.84 2.35 1.22 ;
      LAYER VIA1 ;
        RECT 2.255 1.055 2.345 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.797 1.08 1.192 1.17 ;
      RECT 1.102 0.395 1.192 1.17 ;
      RECT 1.102 0.835 1.825 0.925 ;
      RECT 1.735 0.625 1.825 0.925 ;
      RECT 1.735 0.625 2.075 0.715 ;
      RECT 1.047 0.395 1.192 0.485 ;
      RECT 0.322 0.395 0.912 0.485 ;
      RECT 0.822 0.215 0.912 0.485 ;
      RECT 0.322 0.345 0.412 0.485 ;
      RECT 1.322 0.215 1.412 0.355 ;
      RECT 0.822 0.215 1.412 0.305 ;
  END
END OA22X6H7R

MACRO OA31X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA31X0P5H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.11 1.055 1.2 1.48 ;
        RECT 0.07 1.04 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.085 -0.08 1.225 0.345 ;
        RECT 0.56 -0.08 0.7 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.625 1.035 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.705 0.755 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.625 0.545 0.85 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.39 0.225 1.545 0.375 ;
        RECT 1.39 0.225 1.48 1.16 ;
      LAYER MET2 ;
        RECT 1.45 0.18 1.55 0.56 ;
      LAYER VIA1 ;
        RECT 1.455 0.255 1.545 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.295 1.08 0.945 1.17 ;
      RECT 0.855 0.865 0.945 1.17 ;
      RECT 0.855 0.865 1.3 0.955 ;
      RECT 1.21 0.445 1.3 0.955 ;
      RECT 0.07 0.445 1.3 0.535 ;
      RECT 0.07 0.245 0.16 0.535 ;
      RECT 0.295 0.265 0.965 0.355 ;
  END
END OA31X0P5H7R

MACRO OA31X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA31X0P7H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.115 1.05 1.205 1.48 ;
        RECT 0.075 1.035 0.165 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.09 -0.08 1.23 0.325 ;
        RECT 0.565 -0.08 0.705 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.625 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.75 0.775 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.395 0.625 0.545 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.415 0.225 1.545 0.375 ;
        RECT 1.415 0.225 1.505 1.103 ;
      LAYER MET2 ;
        RECT 1.45 0.18 1.55 0.56 ;
      LAYER VIA1 ;
        RECT 1.455 0.255 1.545 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.3 1.07 1 1.16 ;
      RECT 0.91 0.87 1 1.16 ;
      RECT 0.91 0.87 1.325 0.96 ;
      RECT 1.235 0.445 1.325 0.96 ;
      RECT 0.075 0.445 1.325 0.535 ;
      RECT 0.075 0.225 0.165 0.535 ;
      RECT 0.3 0.265 0.97 0.355 ;
  END
END OA31X0P7H7R

MACRO OA31X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA31X1H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.115 1.05 1.205 1.48 ;
        RECT 0.075 1.035 0.165 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.09 -0.08 1.23 0.345 ;
        RECT 0.565 -0.08 0.705 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.625 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.75 0.775 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.395 0.625 0.545 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.415 0.225 1.545 0.375 ;
        RECT 1.415 0.225 1.505 1.055 ;
      LAYER MET2 ;
        RECT 1.45 0.18 1.55 0.56 ;
      LAYER VIA1 ;
        RECT 1.455 0.255 1.545 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.3 1.07 1 1.16 ;
      RECT 0.91 0.87 1 1.16 ;
      RECT 0.91 0.87 1.325 0.96 ;
      RECT 1.235 0.445 1.325 0.96 ;
      RECT 0.075 0.445 1.325 0.535 ;
      RECT 0.075 0.245 0.165 0.535 ;
      RECT 0.3 0.265 0.97 0.355 ;
  END
END OA31X1H7R

MACRO OA31X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA31X1P4H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.115 1.05 1.205 1.48 ;
        RECT 0.075 1.035 0.165 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.115 -0.08 1.205 0.35 ;
        RECT 0.565 -0.08 0.705 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.625 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.75 0.775 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.395 0.625 0.545 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.415 0.225 1.545 0.375 ;
        RECT 1.415 0.225 1.505 1.011 ;
      LAYER MET2 ;
        RECT 1.45 0.18 1.55 0.56 ;
      LAYER VIA1 ;
        RECT 1.455 0.255 1.545 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.3 1.07 1 1.16 ;
      RECT 0.91 0.87 1 1.16 ;
      RECT 0.91 0.87 1.325 0.96 ;
      RECT 1.235 0.445 1.325 0.96 ;
      RECT 0.075 0.445 1.325 0.535 ;
      RECT 0.075 0.225 0.165 0.535 ;
      RECT 0.3 0.265 0.97 0.355 ;
  END
END OA31X1P4H7R

MACRO OA31X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA31X2H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.615 1.055 1.705 1.48 ;
        RECT 1.1 1.07 1.19 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.605 -0.08 1.745 0.205 ;
        RECT 1.075 -0.08 1.215 0.355 ;
        RECT 0.56 -0.08 0.7 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.625 1.035 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.705 0.755 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.365 0.625 0.545 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.36 0.795 1.745 0.885 ;
        RECT 1.655 0.295 1.745 0.885 ;
        RECT 1.325 0.295 1.745 0.385 ;
        RECT 1.36 0.795 1.45 1.14 ;
      LAYER MET2 ;
        RECT 1.65 0.23 1.75 0.76 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.295 1.07 0.96 1.16 ;
      RECT 0.87 0.885 0.96 1.16 ;
      RECT 0.87 0.885 1.215 0.975 ;
      RECT 1.125 0.445 1.215 0.975 ;
      RECT 1.125 0.535 1.565 0.625 ;
      RECT 0.07 0.445 1.215 0.535 ;
      RECT 0.07 0.255 0.16 0.535 ;
      RECT 0.295 0.265 0.965 0.355 ;
  END
END OA31X2H7R

MACRO OA31X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA31X3H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.6 1.055 1.69 1.48 ;
        RECT 1.1 1.07 1.19 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.59 -0.08 1.73 0.25 ;
        RECT 1.1 -0.08 1.19 0.35 ;
        RECT 0.56 -0.08 0.7 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.625 1.035 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.705 0.755 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.365 0.625 0.545 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.35 0.795 1.745 0.885 ;
        RECT 1.655 0.34 1.745 0.885 ;
        RECT 1.325 0.34 1.745 0.43 ;
        RECT 1.35 0.795 1.44 1.045 ;
      LAYER MET2 ;
        RECT 1.65 0.23 1.75 0.76 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.295 1.07 0.96 1.16 ;
      RECT 0.87 0.885 0.96 1.16 ;
      RECT 0.87 0.885 1.215 0.975 ;
      RECT 1.125 0.445 1.215 0.975 ;
      RECT 1.125 0.615 1.565 0.705 ;
      RECT 0.07 0.445 1.215 0.535 ;
      RECT 0.07 0.255 0.16 0.535 ;
      RECT 0.295 0.265 0.965 0.355 ;
  END
END OA31X3H7R

MACRO OA31X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA31X4H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.615 1.055 1.705 1.48 ;
        RECT 1.1 1.07 1.19 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.575 -0.08 1.715 0.305 ;
        RECT 1.1 -0.08 1.19 0.35 ;
        RECT 0.56 -0.08 0.7 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.625 1.035 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.685 0.755 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.365 0.625 0.545 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.325 0.835 1.745 0.925 ;
        RECT 1.655 0.395 1.745 0.925 ;
        RECT 1.325 0.395 1.745 0.485 ;
      LAYER MET2 ;
        RECT 1.65 0.23 1.75 0.76 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.295 1.07 0.96 1.16 ;
      RECT 0.87 0.885 0.96 1.16 ;
      RECT 0.87 0.885 1.215 0.975 ;
      RECT 1.125 0.445 1.215 0.975 ;
      RECT 1.125 0.625 1.565 0.715 ;
      RECT 0.07 0.445 1.215 0.535 ;
      RECT 0.07 0.305 0.16 0.535 ;
      RECT 0.295 0.265 0.965 0.355 ;
  END
END OA31X4H7R

MACRO OAI211X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211X0P5H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.795 1.05 0.885 1.48 ;
        RECT 0.07 0.87 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.395 0.6 0.545 0.78 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.675 0.655 0.975 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.425 1.145 0.575 ;
        RECT 0.925 0.425 1.145 0.53 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.505 0.87 1.345 0.96 ;
        RECT 1.255 0.225 1.345 0.96 ;
        RECT 1.045 0.225 1.345 0.32 ;
      LAYER MET2 ;
        RECT 1.25 0.18 1.35 0.56 ;
      LAYER VIA1 ;
        RECT 1.255 0.255 1.345 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.42 0.66 0.51 ;
      RECT 0.57 0.22 0.66 0.51 ;
      RECT 0.07 0.205 0.16 0.51 ;
  END
END OAI211X0P5H7R

MACRO OAI211X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211X0P7H7R 0 0 ;
  SIZE 1.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.2 1.48 ;
        RECT 1.005 1.08 1.145 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.2 0.08 ;
        RECT 0.755 -0.08 0.895 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.035 0.75 1.155 0.975 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.7 0.625 0.945 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.435 0.555 0.555 0.78 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.535 0.16 0.795 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.57 0.915 0.66 1.108 ;
        RECT 0.07 0.915 0.66 1.005 ;
        RECT 0.255 0.255 0.345 1.005 ;
        RECT 0.045 0.255 0.345 0.345 ;
        RECT 0.07 0.915 0.16 1.123 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.639 0.395 1.12 0.485 ;
      RECT 1.03 0.23 1.12 0.485 ;
      RECT 0.62 0.347 0.639 0.476 ;
      RECT 0.576 0.395 1.12 0.444 ;
      RECT 0.53 0.235 0.62 0.399 ;
      RECT 0.53 0.376 0.677 0.399 ;
  END
END OAI211X0P7H7R

MACRO OAI211X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211X1H7R 0 0 ;
  SIZE 1.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.2 1.48 ;
        RECT 1.005 1.08 1.145 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.2 0.08 ;
        RECT 0.755 -0.08 0.895 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.035 0.725 1.145 0.975 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.7 0.625 0.945 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.435 0.595 0.555 0.82 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.545 0.165 0.795 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.57 0.915 0.66 1.06 ;
        RECT 0.07 0.915 0.66 1.005 ;
        RECT 0.255 0.29 0.345 1.005 ;
        RECT 0.045 0.29 0.345 0.38 ;
        RECT 0.07 0.915 0.16 1.075 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.53 0.395 1.12 0.485 ;
      RECT 1.03 0.265 1.12 0.485 ;
      RECT 0.53 0.28 0.62 0.485 ;
  END
END OAI211X1H7R

MACRO OAI211X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211X1P4H7R 0 0 ;
  SIZE 1.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.2 1.48 ;
        RECT 1.005 1.08 1.145 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.2 0.08 ;
        RECT 0.755 -0.08 0.895 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.035 0.68 1.145 0.975 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.7 0.625 0.945 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.435 0.6 0.555 0.825 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.535 0.165 0.785 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.07 0.915 0.685 1.005 ;
        RECT 0.255 0.325 0.345 1.005 ;
        RECT 0.045 0.325 0.345 0.415 ;
        RECT 0.07 0.915 0.16 1.058 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.53 0.395 1.12 0.485 ;
      RECT 1.03 0.3 1.12 0.485 ;
      RECT 0.53 0.315 0.62 0.485 ;
  END
END OAI211X1P4H7R

MACRO OAI211X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211X2H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.257 1.08 1.397 1.48 ;
        RECT 0.572 1.07 0.662 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.007 -0.08 1.147 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.64 1.345 0.975 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.952 0.615 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.58 0.79 0.78 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.575 0.385 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.297 0.885 0.937 0.975 ;
        RECT 0.297 0.255 0.575 0.345 ;
        RECT 0.475 0.255 0.565 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.18 0.55 0.56 ;
      LAYER VIA1 ;
        RECT 0.455 0.255 0.545 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.757 0.395 1.372 0.485 ;
      RECT 1.282 0.345 1.372 0.485 ;
  END
END OAI211X2H7R

MACRO OAI211X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211X3H7R 0 0 ;
  SIZE 2.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.8 1.48 ;
        RECT 2.025 1.095 2.165 1.48 ;
        RECT 0.795 1.095 0.935 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.8 0.08 ;
        RECT 2.085 -0.08 2.225 0.305 ;
        RECT 1.585 -0.08 1.725 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.955 0.655 2.295 0.745 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.225 0.655 1.765 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.725 0.655 1.065 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.245 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 1.11 1.685 1.2 ;
        RECT 1.545 1.08 1.685 1.2 ;
        RECT 1.055 0.915 1.16 1.2 ;
        RECT 0.07 0.915 1.16 1.005 ;
        RECT 0.545 0.915 0.685 1.02 ;
        RECT 0.36 0.35 0.45 1.005 ;
        RECT 0.31 0.35 0.45 0.44 ;
        RECT 0.07 0.915 0.16 1.06 ;
      LAYER MET2 ;
        RECT 1.05 0.84 1.15 1.22 ;
      LAYER VIA1 ;
        RECT 1.055 1.055 1.145 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.84 0.455 1.45 0.545 ;
      RECT 1.36 0.28 1.45 0.545 ;
      RECT 2.36 0.28 2.45 0.5 ;
      RECT 1.36 0.41 2.45 0.5 ;
      RECT 0.84 0.35 0.98 0.545 ;
      RECT 1.86 0.295 1.95 0.5 ;
      RECT 2.3 0.9 2.39 1.06 ;
      RECT 1.775 0.9 1.915 1.035 ;
      RECT 1.295 0.9 1.435 1.02 ;
      RECT 1.295 0.9 2.39 0.99 ;
      RECT 0.07 0.17 0.16 0.41 ;
      RECT 0.575 0.17 0.715 0.37 ;
      RECT 1.105 0.17 1.245 0.365 ;
      RECT 0.07 0.17 1.245 0.26 ;
  END
END OAI211X3H7R

MACRO OAI211X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211X4H7R 0 0 ;
  SIZE 3 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3 1.48 ;
        RECT 2.302 1.07 2.392 1.48 ;
        RECT 1.072 1.07 1.162 1.48 ;
        RECT 0.572 1.07 0.662 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3 0.08 ;
        RECT 2.277 -0.08 2.417 0.305 ;
        RECT 1.777 -0.08 1.917 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.207 0.655 2.547 0.745 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.447 0.655 1.987 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.917 0.655 1.257 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.365 0.625 0.545 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.322 1.055 1.937 1.145 ;
        RECT 1.322 0.865 1.412 1.205 ;
        RECT 0.297 0.865 1.412 0.955 ;
        RECT 0.822 0.865 0.912 1.18 ;
        RECT 0.635 0.395 0.725 0.955 ;
        RECT 0.547 0.395 0.725 0.485 ;
        RECT 0.297 0.865 0.412 1.18 ;
      LAYER MET2 ;
        RECT 1.45 0.84 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.047 0.41 2.642 0.5 ;
      RECT 2.552 0.355 2.642 0.5 ;
      RECT 2.027 0.395 2.167 0.5 ;
      RECT 1.552 0.355 1.642 0.5 ;
      RECT 1.047 0.395 1.187 0.5 ;
      RECT 2.552 0.85 2.642 1.19 ;
      RECT 2.052 0.85 2.142 1.165 ;
      RECT 1.547 0.85 1.687 0.955 ;
      RECT 1.547 0.85 2.642 0.94 ;
      RECT 0.322 0.215 0.412 0.355 ;
      RECT 1.297 0.215 1.437 0.32 ;
      RECT 0.322 0.215 1.437 0.305 ;
  END
END OAI211X4H7R

MACRO OAI211X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211X6H7R 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.8 1.48 ;
        RECT 3.322 0.855 3.412 1.48 ;
        RECT 2.822 1.07 2.912 1.48 ;
        RECT 1.572 1.07 1.662 1.48 ;
        RECT 1.072 1.07 1.162 1.48 ;
        RECT 0.572 1.07 0.662 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.8 0.08 ;
        RECT 3.047 -0.08 3.187 0.305 ;
        RECT 2.547 -0.08 2.687 0.305 ;
        RECT 2.047 -0.08 2.187 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.727 0.655 3.267 0.745 ;
      LAYER MET2 ;
        RECT 2.85 0.43 2.95 0.96 ;
      LAYER VIA1 ;
        RECT 2.855 0.655 2.945 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.957 0.655 2.497 0.745 ;
      LAYER MET2 ;
        RECT 2.05 0.255 2.15 0.785 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.227 0.655 1.767 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.502 0.655 1.042 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.822 1.055 2.437 1.145 ;
        RECT 1.822 0.855 1.912 1.195 ;
        RECT 0.322 0.855 1.912 0.945 ;
        RECT 1.322 0.855 1.412 1.2 ;
        RECT 0.322 0.395 0.937 0.485 ;
        RECT 0.822 0.855 0.912 1.195 ;
        RECT 0.322 0.355 0.412 1.165 ;
      LAYER MET2 ;
        RECT 2.05 1.015 2.15 1.22 ;
      LAYER VIA1 ;
        RECT 2.055 1.055 2.145 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.297 0.395 3.412 0.485 ;
      RECT 3.322 0.345 3.412 0.485 ;
      RECT 3.072 0.87 3.162 1.21 ;
      RECT 2.572 0.87 2.662 1.185 ;
      RECT 2.047 0.87 3.162 0.96 ;
      RECT 0.547 0.215 1.687 0.305 ;
  END
END OAI211X6H7R

MACRO OAI21BX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21BX0P5H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.815 1.07 0.905 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.05 -0.08 1.14 0.345 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.61 0.19 0.81 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.775 0.545 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.045 0.55 1.165 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.635 0.525 0.945 0.615 ;
        RECT 0.855 0.23 0.945 0.615 ;
        RECT 0.795 0.23 0.945 0.32 ;
        RECT 0.505 1.065 0.725 1.155 ;
        RECT 0.635 0.525 0.725 1.155 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.145 0.865 1.235 1.155 ;
      RECT 0.815 0.865 1.39 0.955 ;
      RECT 1.3 0.205 1.39 0.955 ;
      RECT 0.815 0.805 0.905 0.955 ;
      RECT 0.07 0.395 0.511 0.485 ;
      RECT 0.07 0.395 0.557 0.462 ;
      RECT 0.473 0.376 0.616 0.403 ;
      RECT 0.557 0.304 0.57 0.433 ;
      RECT 0.07 0.205 0.16 0.485 ;
      RECT 0.511 0.334 0.616 0.403 ;
      RECT 0.57 0.19 0.66 0.358 ;
  END
END OAI21BX0P5H7R

MACRO OAI21BX0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21BX0P7H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.815 1.07 0.905 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.05 -0.08 1.14 0.345 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.61 0.19 0.81 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.415 0.765 0.545 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.55 1.175 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.635 0.505 0.945 0.595 ;
        RECT 0.855 0.255 0.945 0.595 ;
        RECT 0.795 0.255 0.945 0.345 ;
        RECT 0.505 1.065 0.725 1.155 ;
        RECT 0.635 0.505 0.725 1.155 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.145 0.865 1.235 1.155 ;
      RECT 0.815 0.865 1.39 0.955 ;
      RECT 1.3 0.205 1.39 0.955 ;
      RECT 0.815 0.77 0.905 0.955 ;
      RECT 0.07 0.395 0.511 0.485 ;
      RECT 0.07 0.395 0.557 0.462 ;
      RECT 0.473 0.376 0.616 0.403 ;
      RECT 0.557 0.304 0.57 0.433 ;
      RECT 0.07 0.205 0.16 0.485 ;
      RECT 0.511 0.334 0.616 0.403 ;
      RECT 0.57 0.19 0.66 0.358 ;
  END
END OAI21BX0P7H7R

MACRO OAI21BX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21BX1H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.815 1.07 0.905 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.05 -0.08 1.14 0.345 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.61 0.19 0.81 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.705 0.545 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.55 1.175 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.635 0.515 0.945 0.605 ;
        RECT 0.855 0.29 0.945 0.605 ;
        RECT 0.795 0.29 0.945 0.38 ;
        RECT 0.505 1.065 0.725 1.155 ;
        RECT 0.635 0.515 0.725 1.155 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.145 0.865 1.235 1.155 ;
      RECT 0.815 0.865 1.39 0.955 ;
      RECT 1.3 0.205 1.39 0.955 ;
      RECT 0.815 0.725 0.905 0.955 ;
      RECT 0.07 0.395 0.511 0.485 ;
      RECT 0.07 0.395 0.557 0.462 ;
      RECT 0.473 0.376 0.616 0.403 ;
      RECT 0.557 0.304 0.57 0.433 ;
      RECT 0.07 0.265 0.16 0.485 ;
      RECT 0.511 0.334 0.616 0.403 ;
      RECT 0.57 0.19 0.66 0.358 ;
  END
END OAI21BX1H7R

MACRO OAI21BX1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21BX1P4H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.815 1.07 0.905 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.05 -0.08 1.14 0.345 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.68 0.545 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.55 1.175 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.635 0.49 0.945 0.58 ;
        RECT 0.82 0.3 0.945 0.58 ;
        RECT 0.505 1.065 0.725 1.155 ;
        RECT 0.635 0.49 0.725 1.155 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.145 0.865 1.235 1.155 ;
      RECT 0.815 0.865 1.39 0.955 ;
      RECT 1.3 0.205 1.39 0.955 ;
      RECT 0.815 0.68 0.905 0.955 ;
      RECT 0.07 0.395 0.511 0.485 ;
      RECT 0.07 0.395 0.557 0.462 ;
      RECT 0.473 0.376 0.616 0.403 ;
      RECT 0.557 0.304 0.57 0.433 ;
      RECT 0.07 0.205 0.16 0.485 ;
      RECT 0.511 0.334 0.616 0.403 ;
      RECT 0.57 0.19 0.66 0.358 ;
  END
END OAI21BX1P4H7R

MACRO OAI21BX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21BX2H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.067 1.07 1.157 1.48 ;
        RECT 0.322 1.055 0.412 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.302 -0.08 1.392 0.345 ;
        RECT 0.547 -0.08 0.687 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.22 0.655 0.52 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.575 0.775 0.8 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.625 1.435 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.205 1.162 0.37 ;
        RECT 1.055 0.205 1.147 0.4 ;
        RECT 0.977 0.396 1.101 0.446 ;
        RECT 1.023 0.357 1.055 0.485 ;
        RECT 0.933 0.441 1.023 0.524 ;
        RECT 0.757 0.89 0.977 0.98 ;
        RECT 0.887 0.486 0.977 0.98 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.56 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.397 0.865 1.487 1.155 ;
      RECT 1.067 0.865 1.642 0.955 ;
      RECT 1.552 0.205 1.642 0.955 ;
      RECT 1.067 0.61 1.157 0.955 ;
      RECT 0.322 0.395 0.763 0.485 ;
      RECT 0.322 0.395 0.809 0.462 ;
      RECT 0.725 0.376 0.868 0.403 ;
      RECT 0.809 0.304 0.822 0.433 ;
      RECT 0.322 0.345 0.412 0.485 ;
      RECT 0.763 0.334 0.868 0.403 ;
      RECT 0.822 0.19 0.912 0.358 ;
  END
END OAI21BX2H7R

MACRO OAI21BX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21BX3H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 1.83 1.07 1.92 1.48 ;
        RECT 1.24 1.11 1.38 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 2.34 -0.08 2.43 0.345 ;
        RECT 0.99 -0.08 1.13 0.175 ;
        RECT 0.36 -0.08 0.5 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.14 0.455 1.23 0.605 ;
        RECT 0.17 0.455 1.23 0.545 ;
        RECT 0.17 0.455 0.26 0.63 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.475 0.655 0.815 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.112 0.655 2.412 0.745 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.554 0.35 1.71 0.44 ;
        RECT 0.545 0.93 1.695 1.02 ;
        RECT 1.455 0.426 1.592 0.459 ;
        RECT 1.501 0.381 1.71 0.44 ;
        RECT 1.545 0.354 1.554 0.483 ;
        RECT 1.455 0.426 1.545 1.02 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.08 0.89 2.17 1.195 ;
      RECT 1.805 0.89 2.17 0.98 ;
      RECT 1.805 0.666 1.895 0.98 ;
      RECT 1.655 0.7 1.895 0.79 ;
      RECT 1.794 0.694 1.895 0.79 ;
      RECT 1.851 0.621 1.941 0.704 ;
      RECT 1.895 0.576 1.987 0.658 ;
      RECT 1.941 0.53 2.033 0.612 ;
      RECT 1.941 0.53 2.079 0.566 ;
      RECT 1.987 0.484 2.09 0.538 ;
      RECT 2.033 0.438 2.136 0.509 ;
      RECT 2.079 0.409 2.09 0.538 ;
      RECT 2.09 0.205 2.18 0.464 ;
      RECT 0.045 0.265 1.42 0.355 ;
      RECT 1.33 0.17 1.42 0.355 ;
      RECT 1.86 0.17 1.95 0.345 ;
      RECT 1.33 0.17 1.95 0.26 ;
      RECT 0.295 1.11 1 1.2 ;
      RECT 0.295 1.095 0.435 1.2 ;
  END
END OAI21BX3H7R

MACRO OAI21BX4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21BX4H7R 0 0 ;
  SIZE 2.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.8 1.48 ;
        RECT 2.082 1.07 2.172 1.48 ;
        RECT 1.517 1.07 1.607 1.48 ;
        RECT 0.402 1.055 0.492 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.8 0.08 ;
        RECT 2.562 -0.08 2.652 0.345 ;
        RECT 1.242 -0.08 1.382 0.175 ;
        RECT 0.612 -0.08 0.752 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.392 0.455 1.482 0.68 ;
        RECT 0.502 0.455 1.482 0.545 ;
        RECT 0.502 0.455 0.592 0.71 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.797 0.655 1.137 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.357 0.655 2.657 0.745 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.927 0.885 1.947 0.975 ;
        RECT 1.761 0.395 1.947 0.485 ;
        RECT 1.655 0.478 1.799 0.504 ;
        RECT 1.701 0.433 1.947 0.485 ;
        RECT 1.745 0.403 1.761 0.531 ;
        RECT 1.655 0.478 1.745 0.975 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.332 0.89 2.422 1.035 ;
      RECT 2.065 0.89 2.422 0.98 ;
      RECT 2.065 0.655 2.155 0.98 ;
      RECT 1.877 0.655 2.155 0.745 ;
      RECT 2.066 0.632 2.201 0.671 ;
      RECT 2.112 0.587 2.201 0.671 ;
      RECT 2.155 0.543 2.247 0.625 ;
      RECT 2.155 0.543 2.293 0.579 ;
      RECT 2.201 0.497 2.312 0.547 ;
      RECT 2.247 0.451 2.358 0.514 ;
      RECT 2.293 0.418 2.312 0.547 ;
      RECT 2.312 0.305 2.402 0.469 ;
      RECT 0.297 0.265 1.672 0.355 ;
      RECT 1.582 0.17 1.672 0.355 ;
      RECT 2.082 0.17 2.172 0.345 ;
      RECT 1.582 0.17 2.172 0.26 ;
      RECT 0.677 1.095 1.317 1.185 ;
  END
END OAI21BX4H7R

MACRO OAI21BX6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21BX6H7R 0 0 ;
  SIZE 3.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.4 1.48 ;
        RECT 2.535 1.07 2.625 1.48 ;
        RECT 2.035 1.07 2.125 1.48 ;
        RECT 0.785 1.07 0.875 1.48 ;
        RECT 0.285 0.855 0.375 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.4 0.08 ;
        RECT 3.015 -0.08 3.105 0.345 ;
        RECT 1.51 -0.08 1.65 0.305 ;
        RECT 1.01 -0.08 1.15 0.305 ;
        RECT 0.51 -0.08 0.65 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.655 0.98 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.19 0.655 1.73 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.81 0.65 3.045 0.765 ;
      LAYER MET2 ;
        RECT 2.85 0.43 2.95 0.96 ;
      LAYER VIA1 ;
        RECT 2.855 0.655 2.945 0.745 ;
    END
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.535 0.295 2.625 0.437 ;
        RECT 1.95 0.395 2.623 0.461 ;
        RECT 1.95 0.395 2.577 0.485 ;
        RECT 2.285 0.855 2.375 1.195 ;
        RECT 1.285 0.855 2.375 0.945 ;
        RECT 1.95 0.395 2.04 0.945 ;
        RECT 1.785 0.855 1.875 1.195 ;
        RECT 1.285 0.855 1.375 1 ;
      LAYER MET2 ;
        RECT 2.05 0.63 2.15 1.16 ;
      LAYER VIA1 ;
        RECT 2.055 0.855 2.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.785 0.855 2.875 1.195 ;
      RECT 2.575 0.855 2.875 0.945 ;
      RECT 2.575 0.602 2.665 0.945 ;
      RECT 2.13 0.625 2.665 0.715 ;
      RECT 2.621 0.557 2.711 0.64 ;
      RECT 2.621 0.557 2.757 0.594 ;
      RECT 2.665 0.512 2.765 0.567 ;
      RECT 2.711 0.466 2.811 0.54 ;
      RECT 2.757 0.439 2.765 0.567 ;
      RECT 2.765 0.329 2.855 0.495 ;
      RECT 0.285 0.395 1.85 0.485 ;
      RECT 1.76 0.215 1.85 0.485 ;
      RECT 0.285 0.33 0.375 0.485 ;
      RECT 1.76 0.215 2.4 0.305 ;
      RECT 1.035 1.095 1.65 1.185 ;
      RECT 1.035 0.845 1.125 1.185 ;
      RECT 0.51 0.885 1.125 0.975 ;
  END
END OAI21BX6H7R

MACRO OAI21X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X0P5H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.815 1.215 0.955 1.48 ;
        RECT 0.07 0.985 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.295 -0.08 0.435 0.34 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.245 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.38 0.855 0.575 0.945 ;
        RECT 0.38 0.775 0.505 0.945 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.61 0.75 0.81 ;
        RECT 0.575 0.61 0.75 0.715 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.53 1.035 0.945 1.125 ;
        RECT 0.84 0.225 0.945 1.125 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.56 ;
      LAYER VIA1 ;
        RECT 0.855 0.255 0.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.43 0.66 0.52 ;
      RECT 0.57 0.255 0.66 0.52 ;
      RECT 0.07 0.24 0.16 0.52 ;
  END
END OAI21X0P5H7R

MACRO OAI21X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X0P7H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.84 1.115 0.93 1.48 ;
        RECT 0.07 0.985 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.295 -0.08 0.435 0.355 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.245 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.415 0.855 0.575 0.945 ;
        RECT 0.415 0.715 0.505 0.945 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.65 0.625 0.765 0.8 ;
        RECT 0.595 0.625 0.765 0.75 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.305 0.945 0.901 ;
        RECT 0.745 0.928 0.855 0.978 ;
        RECT 0.791 0.882 0.901 0.946 ;
        RECT 0.837 0.85 0.855 0.978 ;
        RECT 0.795 0.305 0.945 0.395 ;
        RECT 0.699 0.974 0.837 1.01 ;
        RECT 0.661 1.016 0.791 1.056 ;
        RECT 0.699 0.974 0.791 1.056 ;
        RECT 0.53 1.035 0.745 1.102 ;
        RECT 0.53 1.035 0.699 1.125 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.445 0.66 0.535 ;
      RECT 0.57 0.295 0.66 0.535 ;
      RECT 0.07 0.28 0.16 0.535 ;
  END
END OAI21X0P7H7R

MACRO OAI21X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X1H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.795 1.09 0.935 1.48 ;
        RECT 0.07 1.05 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.26 0.745 ;
        RECT 0.055 0.625 0.145 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 0.72 0.49 0.88 ;
        RECT 0.225 0.855 0.451 0.922 ;
        RECT 0.225 0.855 0.405 0.945 ;
        RECT 0.367 0.838 0.49 0.88 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.595 0.595 0.745 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.57 0.905 0.945 0.995 ;
        RECT 0.84 0.265 0.945 0.995 ;
        RECT 0.57 0.905 0.66 1.055 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.395 0.66 0.485 ;
      RECT 0.57 0.28 0.66 0.485 ;
      RECT 0.07 0.265 0.16 0.485 ;
  END
END OAI21X1H7R

MACRO OAI21X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X1P4H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.795 1.095 0.935 1.48 ;
        RECT 0.07 1.05 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.295 0.715 ;
        RECT 0.055 0.625 0.145 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 0.681 0.49 0.88 ;
        RECT 0.225 0.855 0.451 0.922 ;
        RECT 0.225 0.855 0.405 0.945 ;
        RECT 0.367 0.838 0.49 0.88 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.595 0.595 0.745 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.57 0.905 0.945 0.995 ;
        RECT 0.84 0.3 0.945 0.995 ;
        RECT 0.57 0.905 0.66 1.06 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.395 0.66 0.485 ;
      RECT 0.57 0.315 0.66 0.485 ;
      RECT 0.07 0.3 0.16 0.485 ;
  END
END OAI21X1P4H7R

MACRO OAI21X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X2H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.05 1.095 1.19 1.48 ;
        RECT 0.325 1.05 0.415 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.55 -0.08 0.69 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.655 0.525 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.615 0.745 0.807 ;
        RECT 0.547 0.836 0.655 0.887 ;
        RECT 0.585 0.794 0.701 0.852 ;
        RECT 0.631 0.759 0.655 0.887 ;
        RECT 0.425 0.855 0.631 0.922 ;
        RECT 0.425 0.855 0.585 0.945 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.85 0.595 1 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.25 0.95 0.785 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.915 1.185 1.005 ;
        RECT 1.095 0.355 1.185 1.005 ;
        RECT 0.825 0.915 0.945 1.175 ;
      LAYER MET2 ;
        RECT 0.85 1.015 0.95 1.22 ;
      LAYER VIA1 ;
        RECT 0.855 1.055 0.945 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.325 0.395 0.94 0.485 ;
      RECT 0.325 0.345 0.415 0.485 ;
  END
END OAI21X2H7R

MACRO OAI21X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X3H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.8 1.055 1.89 1.48 ;
        RECT 1.275 1.08 1.415 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 0.795 -0.08 0.935 0.305 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.195 0.655 0.535 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.695 0.655 1.035 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.435 0.655 1.775 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.55 0.9 1.64 1.045 ;
        RECT 0.795 0.9 1.64 0.99 ;
        RECT 1.255 0.35 1.465 0.44 ;
        RECT 1.255 0.35 1.345 0.99 ;
        RECT 0.795 0.9 0.935 1.02 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.395 1.16 0.485 ;
      RECT 1.07 0.17 1.16 0.485 ;
      RECT 0.57 0.295 0.66 0.485 ;
      RECT 0.07 0.28 0.16 0.485 ;
      RECT 1.63 0.17 1.72 0.345 ;
      RECT 1.07 0.17 1.72 0.26 ;
      RECT 0.57 1.11 1.185 1.2 ;
      RECT 1.045 1.08 1.185 1.2 ;
      RECT 0.57 0.905 0.66 1.2 ;
      RECT 0.07 0.905 0.16 1.06 ;
      RECT 0.07 0.905 0.66 0.995 ;
  END
END OAI21X3H7R

MACRO OAI21X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X4H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 2.052 1.055 2.142 1.48 ;
        RECT 1.552 1.055 1.642 1.48 ;
        RECT 0.547 1.095 0.687 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 1.047 -0.08 1.187 0.305 ;
        RECT 0.547 -0.08 0.687 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.447 0.64 0.787 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.947 0.64 1.287 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.835 0.575 1.97 0.775 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.047 0.865 1.917 0.955 ;
        RECT 1.655 0.35 1.745 0.955 ;
        RECT 1.577 0.35 1.745 0.44 ;
      LAYER MET2 ;
        RECT 1.65 0.23 1.75 0.76 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.322 0.395 1.412 0.485 ;
      RECT 1.322 0.17 1.412 0.485 ;
      RECT 0.322 0.345 0.412 0.485 ;
      RECT 1.882 0.17 1.972 0.345 ;
      RECT 1.322 0.17 1.972 0.26 ;
      RECT 0.822 1.045 1.437 1.135 ;
      RECT 0.822 0.905 0.912 1.135 ;
      RECT 0.297 0.905 0.912 0.995 ;
  END
END OAI21X4H7R

MACRO OAI21X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X6H7R 0 0 ;
  SIZE 3 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3 1.48 ;
        RECT 2.572 0.855 2.662 1.48 ;
        RECT 2.072 1.07 2.162 1.48 ;
        RECT 0.797 1.095 0.937 1.48 ;
        RECT 0.322 0.855 0.412 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3 0.08 ;
        RECT 1.547 -0.08 1.687 0.305 ;
        RECT 1.047 -0.08 1.187 0.305 ;
        RECT 0.547 -0.08 0.687 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.477 0.655 1.017 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.227 0.655 1.767 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.365 0.635 2.59 0.755 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.047 0.395 2.687 0.485 ;
        RECT 2.547 0.38 2.687 0.485 ;
        RECT 1.297 0.885 2.437 0.975 ;
        RECT 2.055 0.395 2.145 0.975 ;
      LAYER MET2 ;
        RECT 2.05 0.63 2.15 1.16 ;
      LAYER VIA1 ;
        RECT 2.055 0.855 2.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.322 0.395 1.912 0.485 ;
      RECT 1.822 0.215 1.912 0.485 ;
      RECT 0.322 0.345 0.412 0.485 ;
      RECT 1.822 0.215 2.437 0.305 ;
      RECT 1.072 1.08 1.687 1.17 ;
      RECT 1.072 0.905 1.162 1.17 ;
      RECT 0.547 0.905 1.162 0.995 ;
  END
END OAI21X6H7R

MACRO OAI21X8H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X8H7R 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.8 1.48 ;
        RECT 3.552 0.855 3.642 1.48 ;
        RECT 3.052 1.07 3.142 1.48 ;
        RECT 2.527 1.08 2.667 1.48 ;
        RECT 1.072 1.07 1.162 1.48 ;
        RECT 0.572 1.07 0.662 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.8 0.08 ;
        RECT 2.047 -0.08 2.187 0.305 ;
        RECT 1.547 -0.08 1.687 0.305 ;
        RECT 1.047 -0.08 1.187 0.305 ;
        RECT 0.547 -0.08 0.687 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.517 0.655 1.257 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.477 0.655 2.217 0.745 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.747 0.655 3.487 0.745 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.547 0.885 3.417 0.975 ;
        RECT 2.477 0.395 3.187 0.485 ;
        RECT 2.455 0.825 2.567 0.975 ;
        RECT 2.477 0.395 2.567 0.975 ;
      LAYER MET2 ;
        RECT 2.45 0.625 2.55 1.16 ;
      LAYER VIA1 ;
        RECT 2.455 0.855 2.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.322 0.395 2.387 0.485 ;
      RECT 2.297 0.215 2.387 0.485 ;
      RECT 0.322 0.345 0.412 0.485 ;
      RECT 3.297 0.215 3.437 0.32 ;
      RECT 2.297 0.215 3.437 0.305 ;
      RECT 1.322 1.08 2.437 1.17 ;
      RECT 1.322 0.89 1.412 1.17 ;
      RECT 0.297 0.89 1.412 0.98 ;
  END
END OAI21X8H7R

MACRO OAI221X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221X0P5H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.16 1.225 1.3 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 0.565 -0.08 0.705 0.175 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.75 0.545 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.75 0.825 0.975 0.945 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.09 0.855 1.375 0.945 ;
        RECT 1.09 0.805 1.18 0.945 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.425 0.55 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.605 1.55 1.135 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.615 1.035 1.725 1.125 ;
        RECT 1.635 0.23 1.725 1.125 ;
        RECT 1.425 0.23 1.725 0.345 ;
      LAYER MET2 ;
        RECT 1.45 0.18 1.55 0.385 ;
      LAYER VIA1 ;
        RECT 1.455 0.255 1.545 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.6 0.495 1.29 0.585 ;
      RECT 1.2 0.205 1.29 0.585 ;
      RECT 0.3 0.265 1.025 0.355 ;
  END
END OAI221X0P5H7R

MACRO OAI221X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221X0P7H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.58 1.055 1.67 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.58 -0.08 1.67 0.345 ;
        RECT 1.055 -0.08 1.195 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.855 1.24 0.945 ;
        RECT 1.15 0.77 1.24 0.945 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.41 0.59 1.545 0.79 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.705 0.645 0.975 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.25 0.95 0.785 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.59 0.585 0.79 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.425 0.345 0.65 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 1.055 1.165 1.145 ;
        RECT 0.655 0.915 0.745 1.145 ;
        RECT 0.045 0.915 0.745 1.005 ;
        RECT 0.045 0.915 0.185 1.098 ;
        RECT 0.045 0.25 0.185 0.34 ;
        RECT 0.045 0.25 0.135 1.098 ;
      LAYER MET2 ;
        RECT 0.85 1.015 0.95 1.22 ;
      LAYER VIA1 ;
        RECT 0.855 1.055 0.945 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.56 0.41 1.42 0.5 ;
      RECT 1.33 0.245 1.42 0.5 ;
      RECT 0.56 0.35 0.7 0.5 ;
      RECT 0.32 0.17 0.41 0.33 ;
      RECT 0.825 0.17 0.965 0.32 ;
      RECT 0.32 0.17 0.965 0.26 ;
  END
END OAI221X0P7H7R

MACRO OAI221X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221X1H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.26 1.045 1.4 1.48 ;
        RECT 0.07 0.925 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 0.57 -0.08 0.71 0.26 ;
        RECT 0.07 -0.08 0.16 0.39 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.62 0.545 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.62 0.23 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.62 0.835 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.62 1.285 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.425 0.565 1.575 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.855 1.755 0.945 ;
        RECT 1.665 0.335 1.755 0.945 ;
        RECT 1.575 0.335 1.755 0.425 ;
        RECT 0.57 1.065 1.115 1.155 ;
        RECT 1.025 0.855 1.115 1.155 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.34 0.17 1.43 0.375 ;
      RECT 0.8 0.17 1.43 0.26 ;
      RECT 0.295 0.35 1.205 0.44 ;
  END
END OAI221X1H7R

MACRO OAI221X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221X1P4H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.58 1.055 1.67 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.58 -0.08 1.67 0.345 ;
        RECT 1.055 -0.08 1.195 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.02 0.855 1.24 0.945 ;
        RECT 1.15 0.705 1.24 0.945 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.41 0.59 1.545 0.79 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.725 0.645 0.995 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.59 0.585 0.79 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.425 0.345 0.65 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.525 1.055 1.165 1.145 ;
        RECT 0.525 0.915 0.615 1.145 ;
        RECT 0.045 0.915 0.615 1.005 ;
        RECT 0.045 0.915 0.185 1.006 ;
        RECT 0.045 0.25 0.185 0.34 ;
        RECT 0.045 0.25 0.135 1.006 ;
      LAYER MET2 ;
        RECT 0.65 0.84 0.75 1.22 ;
      LAYER VIA1 ;
        RECT 0.655 1.055 0.745 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.56 0.41 1.42 0.5 ;
      RECT 1.33 0.315 1.42 0.5 ;
      RECT 0.56 0.355 0.7 0.5 ;
      RECT 0.32 0.17 0.41 0.33 ;
      RECT 0.825 0.17 0.965 0.32 ;
      RECT 0.32 0.17 0.965 0.26 ;
  END
END OAI221X1P4H7R

MACRO OAI221X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221X2H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.832 1.055 1.922 1.48 ;
        RECT 0.572 1.07 0.662 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.802 -0.08 1.892 0.345 ;
        RECT 1.277 -0.08 1.417 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.395 0.595 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.675 0.655 1.975 0.745 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.995 0.595 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.595 0.805 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.425 0.545 0.725 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.077 0.865 1.417 1.155 ;
        RECT 0.255 0.865 1.417 0.955 ;
        RECT 0.255 0.245 0.437 0.335 ;
        RECT 0.255 0.245 0.345 0.955 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.797 0.41 1.642 0.5 ;
      RECT 1.552 0.36 1.642 0.5 ;
      RECT 0.797 0.395 0.937 0.5 ;
      RECT 1.047 0.215 1.187 0.32 ;
      RECT 0.547 0.215 1.187 0.305 ;
  END
END OAI221X2H7R

MACRO OAI221X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221X3H7R 0 0 ;
  SIZE 3.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.4 1.48 ;
        RECT 2.94 1.07 3.03 1.48 ;
        RECT 0.57 0.96 1.315 1.05 ;
        RECT 0.57 0.96 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.4 0.08 ;
        RECT 2.845 -0.08 2.985 0.305 ;
        RECT 2.345 -0.08 2.485 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.275 0.655 2.615 0.745 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.775 0.655 3.115 0.745 ;
      LAYER MET2 ;
        RECT 2.85 0.43 2.95 0.96 ;
      LAYER VIA1 ;
        RECT 2.855 0.655 2.945 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.285 0.6 1.825 0.69 ;
        RECT 1.625 0.6 1.775 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.6 1.065 0.69 ;
        RECT 0.655 0.425 0.745 0.69 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.05 0.625 0.23 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.44 0.855 2.53 1.045 ;
        RECT 1.405 0.855 2.53 0.945 ;
        RECT 1.71 0.855 1.8 1.05 ;
        RECT 0.32 0.78 1.495 0.87 ;
        RECT 0.31 0.35 0.45 0.44 ;
        RECT 0.32 0.35 0.41 1.045 ;
      LAYER MET2 ;
        RECT 1.85 0.625 1.95 1.16 ;
      LAYER VIA1 ;
        RECT 1.855 0.855 1.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.19 1.14 2.78 1.23 ;
      RECT 2.69 0.89 2.78 1.23 ;
      RECT 2.19 1.055 2.28 1.23 ;
      RECT 3.19 0.89 3.28 1.06 ;
      RECT 2.69 0.89 3.28 0.98 ;
      RECT 0.84 0.42 3.21 0.51 ;
      RECT 3.12 0.28 3.21 0.51 ;
      RECT 2.12 0.41 3.21 0.51 ;
      RECT 1.37 0.35 1.51 0.51 ;
      RECT 0.84 0.35 0.98 0.51 ;
      RECT 2.62 0.295 2.71 0.51 ;
      RECT 2.12 0.28 2.21 0.51 ;
      RECT 0.86 1.14 2.05 1.23 ;
      RECT 1.96 1.055 2.05 1.23 ;
      RECT 1.46 1.055 1.55 1.23 ;
      RECT 0.07 0.17 0.16 0.375 ;
      RECT 1.635 0.17 1.775 0.33 ;
      RECT 1.105 0.17 1.245 0.33 ;
      RECT 0.575 0.17 0.715 0.33 ;
      RECT 0.07 0.17 1.775 0.26 ;
  END
END OAI221X3H7R

MACRO OAI221X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221X4H7R 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.8 1.48 ;
        RECT 3.122 1.055 3.212 1.48 ;
        RECT 0.752 0.96 1.497 1.05 ;
        RECT 0.752 0.96 0.842 1.48 ;
        RECT 0.252 1.055 0.342 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.8 0.08 ;
        RECT 3.027 -0.08 3.167 0.305 ;
        RECT 2.527 -0.08 2.667 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.457 0.655 2.797 0.745 ;
      LAYER MET2 ;
        RECT 2.65 0.43 2.75 0.96 ;
      LAYER VIA1 ;
        RECT 2.655 0.655 2.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.957 0.655 3.297 0.745 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.537 0.59 2.077 0.68 ;
        RECT 1.825 0.59 1.975 0.745 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.59 1.247 0.68 ;
        RECT 0.855 0.425 0.945 0.68 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.232 0.625 0.412 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.597 0.855 2.737 0.975 ;
        RECT 1.587 0.855 2.737 0.945 ;
        RECT 0.502 0.78 1.677 0.87 ;
        RECT 0.502 0.395 0.687 0.485 ;
        RECT 0.502 0.395 0.592 0.95 ;
      LAYER MET2 ;
        RECT 2.05 0.63 2.15 1.16 ;
      LAYER VIA1 ;
        RECT 2.055 0.855 2.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.347 1.065 2.962 1.155 ;
      RECT 2.872 0.875 2.962 1.155 ;
      RECT 2.872 0.875 3.487 0.965 ;
      RECT 1.107 0.41 3.392 0.5 ;
      RECT 3.302 0.355 3.392 0.5 ;
      RECT 2.777 0.395 2.917 0.5 ;
      RECT 2.302 0.355 2.392 0.5 ;
      RECT 1.607 0.36 1.747 0.5 ;
      RECT 1.107 0.36 1.247 0.5 ;
      RECT 1.042 1.14 1.705 1.23 ;
      RECT 1.617 1.08 2.257 1.17 ;
      RECT 0.322 0.18 0.412 0.355 ;
      RECT 1.857 0.18 1.997 0.32 ;
      RECT 1.357 0.18 1.497 0.305 ;
      RECT 0.857 0.18 0.997 0.305 ;
      RECT 0.322 0.18 1.997 0.27 ;
  END
END OAI221X4H7R

MACRO OAI222X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222X0P5H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 2.04 0.925 2.13 1.48 ;
        RECT 1.135 1.115 1.275 1.48 ;
        RECT 0.07 0.925 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 0.35 -0.08 0.44 0.26 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.53 0.555 0.8 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.165 0.625 1.345 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.765 0.625 0.945 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.855 0.675 1.945 0.975 ;
      LAYER MET2 ;
        RECT 1.85 0.625 1.95 1.16 ;
      LAYER VIA1 ;
        RECT 1.855 0.855 1.945 0.945 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.655 0.55 1.745 0.785 ;
        RECT 1.625 0.55 1.745 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.435 0.35 2.105 0.44 ;
        RECT 0.59 0.935 1.545 1.025 ;
        RECT 1.435 0.825 1.545 1.025 ;
        RECT 1.435 0.35 1.525 1.025 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.855 0.17 1.84 0.26 ;
      RECT 0.06 0.35 1.26 0.44 ;
  END
END OAI222X0P5H7R

MACRO OAI222X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222X0P7H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.875 1.055 1.965 1.48 ;
        RECT 1.105 1.225 1.245 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.875 -0.08 1.965 0.345 ;
        RECT 1.35 -0.08 1.49 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.8 0.625 2.015 0.775 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.41 0.795 1.59 0.945 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.82 1.225 0.955 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.685 0.655 0.975 0.745 ;
        RECT 0.685 0.655 0.935 0.765 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.505 0.855 0.775 0.945 ;
        RECT 0.505 0.77 0.595 0.945 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 1.045 1.49 1.135 ;
        RECT 0.325 1.055 0.605 1.145 ;
        RECT 0.31 0.35 0.45 0.44 ;
        RECT 0.325 0.35 0.415 1.145 ;
      LAYER MET2 ;
        RECT 0.45 0.84 0.55 1.22 ;
      LAYER VIA1 ;
        RECT 0.455 1.055 0.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.84 0.475 1.715 0.565 ;
      RECT 1.625 0.245 1.715 0.565 ;
      RECT 0.84 0.35 0.98 0.565 ;
      RECT 0.07 0.17 0.16 0.425 ;
      RECT 0.6 0.17 0.69 0.41 ;
      RECT 1.105 0.17 1.245 0.385 ;
      RECT 0.07 0.17 1.245 0.26 ;
  END
END OAI222X0P7H7R

MACRO OAI222X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222X1H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.99 1.005 2.08 1.48 ;
        RECT 1.16 1.13 1.25 1.48 ;
        RECT 0.07 1.005 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 0.35 -0.08 0.44 0.26 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.53 0.555 0.8 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.165 0.625 1.345 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.765 0.625 0.945 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.965 0.625 2.145 0.775 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.635 0.625 1.875 0.81 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.965 0.35 2.105 0.44 ;
        RECT 1.455 0.445 2.055 0.535 ;
        RECT 1.965 0.35 2.055 0.535 ;
        RECT 1.455 0.35 1.57 0.535 ;
        RECT 0.59 0.91 1.545 1 ;
        RECT 1.455 0.35 1.545 1 ;
        RECT 1.43 0.35 1.57 0.44 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.7 0.17 1.84 0.35 ;
      RECT 0.855 0.17 0.995 0.35 ;
      RECT 0.855 0.17 1.84 0.26 ;
      RECT 0.645 0.445 1.21 0.535 ;
      RECT 1.12 0.35 1.21 0.535 ;
      RECT 0.645 0.35 0.735 0.535 ;
      RECT 1.12 0.35 1.26 0.44 ;
      RECT 0.06 0.35 0.735 0.44 ;
  END
END OAI222X1H7R

MACRO OAI222X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222X1P4H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.86 1.055 1.95 1.48 ;
        RECT 1.105 1.225 1.245 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.86 -0.08 1.95 0.345 ;
        RECT 1.335 -0.08 1.475 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.765 0.625 1.945 0.775 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.425 0.615 1.575 0.795 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.855 1.175 0.945 ;
        RECT 1.035 0.73 1.175 0.945 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.625 0.945 0.775 ;
        RECT 0.735 0.625 0.945 0.765 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.505 0.855 0.775 0.945 ;
        RECT 0.505 0.68 0.595 0.945 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.56 1.045 1.475 1.135 ;
        RECT 0.325 1.055 0.605 1.145 ;
        RECT 0.31 0.35 0.45 0.44 ;
        RECT 0.325 0.35 0.415 1.145 ;
      LAYER MET2 ;
        RECT 0.45 0.84 0.55 1.22 ;
      LAYER VIA1 ;
        RECT 0.455 1.055 0.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.84 0.42 1.7 0.51 ;
      RECT 1.61 0.315 1.7 0.51 ;
      RECT 0.84 0.35 0.98 0.51 ;
      RECT 0.07 0.17 0.16 0.355 ;
      RECT 0.6 0.17 0.69 0.34 ;
      RECT 1.105 0.17 1.245 0.33 ;
      RECT 0.07 0.17 1.245 0.26 ;
  END
END OAI222X1P4H7R

MACRO OAI222X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222X2H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 2.077 1.055 2.167 1.48 ;
        RECT 1.322 1.225 1.462 1.48 ;
        RECT 0.322 1.055 0.412 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 2.052 -0.08 2.142 0.345 ;
        RECT 1.527 -0.08 1.667 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.965 0.625 2.145 0.775 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.655 0.59 1.79 0.79 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.225 0.855 1.375 0.945 ;
        RECT 1.235 0.64 1.325 0.945 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.942 0.615 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.58 0.385 0.78 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.575 0.79 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.749 1.045 1.692 1.135 ;
        RECT 0.766 1.045 0.975 1.145 ;
        RECT 0.657 1.031 0.794 1.059 ;
        RECT 0.657 1.008 0.766 1.059 ;
        RECT 0.749 1.045 0.975 1.137 ;
        RECT 0.611 0.977 0.749 1.013 ;
        RECT 0.703 1.045 1.692 1.105 ;
        RECT 0.611 0.931 0.703 1.013 ;
        RECT 0.541 0.395 0.687 0.485 ;
        RECT 0.541 0.885 0.657 0.932 ;
        RECT 0.521 0.839 0.611 0.91 ;
        RECT 0.565 0.931 0.703 0.967 ;
        RECT 0.475 0.438 0.579 0.492 ;
        RECT 0.475 0.438 0.565 0.877 ;
        RECT 0.521 0.405 0.687 0.485 ;
      LAYER MET2 ;
        RECT 0.85 0.84 0.95 1.22 ;
      LAYER VIA1 ;
        RECT 0.855 1.055 0.945 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.047 0.41 1.892 0.5 ;
      RECT 1.802 0.36 1.892 0.5 ;
      RECT 1.047 0.395 1.187 0.5 ;
      RECT 0.322 0.215 0.412 0.355 ;
      RECT 1.297 0.215 1.437 0.32 ;
      RECT 0.322 0.215 1.437 0.305 ;
  END
END OAI222X2H7R

MACRO OAI222X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222X3H7R 0 0 ;
  SIZE 4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4 1.48 ;
        RECT 3.41 1.055 3.5 1.48 ;
        RECT 2.09 1.225 2.23 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4 0.08 ;
        RECT 3.315 -0.08 3.455 0.305 ;
        RECT 2.815 -0.08 2.955 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.245 0.655 3.585 0.745 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.745 0.655 3.085 0.745 ;
      LAYER MET2 ;
        RECT 2.85 0.43 2.95 0.96 ;
      LAYER VIA1 ;
        RECT 2.855 0.655 2.945 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.955 0.655 2.295 0.745 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.655 1.795 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.655 0.565 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.725 0.655 1.065 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.91 0.865 3 1.05 ;
        RECT 1.55 0.865 3 0.955 ;
        RECT 1.55 0.865 1.64 1.05 ;
        RECT 0.795 0.9 1.64 0.99 ;
        RECT 1.255 0.425 1.345 0.99 ;
        RECT 0.35 0.425 1.345 0.515 ;
        RECT 0.88 0.35 1.02 0.515 ;
        RECT 0.795 0.9 0.935 1.02 ;
        RECT 0.35 0.35 0.49 0.515 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.66 1.14 3.25 1.23 ;
      RECT 3.16 0.875 3.25 1.23 ;
      RECT 2.66 1.055 2.75 1.23 ;
      RECT 3.66 0.875 3.75 1.06 ;
      RECT 3.16 0.875 3.75 0.965 ;
      RECT 1.54 0.44 3.68 0.53 ;
      RECT 3.59 0.28 3.68 0.53 ;
      RECT 3.09 0.295 3.18 0.53 ;
      RECT 2.59 0.28 2.68 0.53 ;
      RECT 2.07 0.35 2.21 0.53 ;
      RECT 1.54 0.35 1.68 0.53 ;
      RECT 1.275 1.14 1.89 1.23 ;
      RECT 1.8 1.045 1.89 1.23 ;
      RECT 2.43 1.045 2.52 1.19 ;
      RECT 1.275 1.08 1.415 1.23 ;
      RECT 1.8 1.045 2.52 1.135 ;
      RECT 0.11 0.17 0.2 0.375 ;
      RECT 2.335 0.17 2.475 0.35 ;
      RECT 1.805 0.17 1.945 0.335 ;
      RECT 1.215 0.17 1.355 0.335 ;
      RECT 0.615 0.17 0.755 0.335 ;
      RECT 0.11 0.17 2.475 0.26 ;
      RECT 0.57 1.11 1.185 1.2 ;
      RECT 1.045 1.08 1.185 1.2 ;
      RECT 0.57 0.915 0.66 1.2 ;
      RECT 0.07 0.915 0.16 1.06 ;
      RECT 0.07 0.915 0.66 1.005 ;
  END
END OAI222X3H7R

MACRO OAI222X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222X4H7R 0 0 ;
  SIZE 4.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.2 1.48 ;
        RECT 3.622 1.055 3.712 1.48 ;
        RECT 2.302 1.225 2.442 1.48 ;
        RECT 0.507 1.095 0.647 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.2 0.08 ;
        RECT 3.527 -0.08 3.667 0.305 ;
        RECT 3.027 -0.08 3.167 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.457 0.655 3.797 0.745 ;
      LAYER MET2 ;
        RECT 3.65 0.43 3.75 0.96 ;
      LAYER VIA1 ;
        RECT 3.655 0.655 3.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.957 0.655 3.297 0.745 ;
      LAYER MET2 ;
        RECT 3.05 0.43 3.15 0.96 ;
      LAYER VIA1 ;
        RECT 3.055 0.655 3.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.167 0.655 2.507 0.745 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.637 0.655 1.977 0.745 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.437 0.655 0.777 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.937 0.655 1.277 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.097 0.855 3.237 0.975 ;
        RECT 1.007 0.855 3.237 0.955 ;
        RECT 1.367 0.395 1.457 0.955 ;
        RECT 0.562 0.395 1.457 0.485 ;
        RECT 1.007 0.855 1.147 0.975 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.847 1.065 3.462 1.155 ;
      RECT 3.372 0.875 3.462 1.155 ;
      RECT 3.372 0.875 3.987 0.965 ;
      RECT 1.752 0.41 3.892 0.5 ;
      RECT 3.802 0.31 3.892 0.5 ;
      RECT 3.277 0.395 3.417 0.5 ;
      RECT 2.802 0.355 2.892 0.5 ;
      RECT 2.282 0.395 2.422 0.5 ;
      RECT 1.752 0.395 1.892 0.5 ;
      RECT 0.322 0.215 0.412 0.355 ;
      RECT 2.547 0.215 2.687 0.32 ;
      RECT 0.322 0.215 2.687 0.305 ;
      RECT 0.782 1.08 1.397 1.17 ;
      RECT 0.782 0.915 0.872 1.17 ;
      RECT 0.257 0.915 0.872 1.005 ;
      RECT 1.487 1.045 2.757 1.135 ;
  END
END OAI222X4H7R

MACRO OAI22X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22X0P5H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.12 1.07 1.21 1.48 ;
        RECT 0.045 1.08 0.185 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.295 -0.08 0.435 0.41 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.825 0.235 0.975 ;
      LAYER MET2 ;
        RECT 0.05 0.625 0.15 1.16 ;
      LAYER VIA1 ;
        RECT 0.055 0.855 0.145 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.75 0.545 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.035 0.75 1.155 0.975 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.64 0.625 0.76 0.85 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.545 1.065 0.945 1.155 ;
        RECT 0.855 0.35 0.945 1.155 ;
        RECT 0.795 0.35 0.945 0.44 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.5 0.514 0.59 ;
      RECT 0.07 0.5 0.56 0.567 ;
      RECT 0.476 0.481 0.616 0.511 ;
      RECT 0.56 0.411 0.57 0.539 ;
      RECT 0.07 0.31 0.16 0.59 ;
      RECT 0.514 0.439 0.616 0.511 ;
      RECT 0.57 0.17 0.66 0.466 ;
      RECT 1.12 0.17 1.21 0.45 ;
      RECT 0.57 0.17 1.21 0.26 ;
  END
END OAI22X0P5H7R

MACRO OAI22X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22X0P7H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.12 1.055 1.21 1.48 ;
        RECT 0.045 1.08 0.185 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.295 -0.08 0.435 0.385 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.75 0.235 0.975 ;
      LAYER MET2 ;
        RECT 0.05 0.625 0.15 1.16 ;
      LAYER VIA1 ;
        RECT 0.055 0.855 0.145 0.945 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.655 0.575 0.755 ;
        RECT 0.425 0.655 0.55 0.905 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.035 0.595 1.155 0.82 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.82 0.76 0.975 ;
        RECT 0.67 0.69 0.76 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.35 0.965 0.44 ;
        RECT 0.545 1.065 0.945 1.155 ;
        RECT 0.855 0.35 0.945 1.155 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.475 0.66 0.565 ;
      RECT 0.57 0.17 0.66 0.565 ;
      RECT 0.07 0.3 0.16 0.565 ;
      RECT 1.13 0.17 1.22 0.425 ;
      RECT 0.57 0.17 1.22 0.26 ;
  END
END OAI22X0P7H7R

MACRO OAI22X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22X1H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.09 1.055 1.18 1.48 ;
        RECT 0.08 1.055 0.17 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.305 -0.08 0.445 0.35 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.705 0.545 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.035 0.625 1.155 0.85 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.645 0.625 0.765 0.85 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 1.065 0.945 1.155 ;
        RECT 0.855 0.35 0.945 1.155 ;
        RECT 0.805 0.35 0.945 0.44 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.08 0.44 0.67 0.53 ;
      RECT 0.58 0.17 0.67 0.53 ;
      RECT 0.08 0.31 0.17 0.53 ;
      RECT 1.09 0.17 1.18 0.39 ;
      RECT 0.58 0.17 1.18 0.26 ;
  END
END OAI22X1H7R

MACRO OAI22X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22X1P4H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.12 1.055 1.21 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.295 -0.08 0.435 0.325 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.395 0.62 0.545 0.855 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.035 0.595 1.155 0.82 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.675 0.745 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.35 0.965 0.44 ;
        RECT 0.545 1.065 0.945 1.155 ;
        RECT 0.855 0.35 0.945 1.155 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.44 0.66 0.53 ;
      RECT 0.57 0.17 0.66 0.53 ;
      RECT 0.07 0.3 0.16 0.53 ;
      RECT 1.13 0.17 1.22 0.385 ;
      RECT 0.57 0.17 1.22 0.26 ;
  END
END OAI22X1P4H7R

MACRO OAI22X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22X2H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.282 1.055 1.372 1.48 ;
        RECT 0.322 1.055 0.412 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 0.547 -0.08 0.687 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.595 0.545 0.795 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.615 0.745 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.282 0.655 1.575 0.745 ;
        RECT 1.282 0.605 1.372 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.615 1.005 0.795 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.757 1.07 1.187 1.16 ;
        RECT 1.097 0.395 1.187 1.16 ;
        RECT 0.915 1.055 1.187 1.16 ;
        RECT 1.047 0.395 1.187 0.485 ;
      LAYER MET2 ;
        RECT 1.05 0.84 1.15 1.22 ;
      LAYER VIA1 ;
        RECT 1.055 1.055 1.145 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.322 0.395 0.912 0.485 ;
      RECT 0.822 0.205 0.912 0.485 ;
      RECT 0.322 0.345 0.412 0.485 ;
      RECT 1.322 0.205 1.412 0.345 ;
      RECT 0.822 0.205 1.412 0.295 ;
  END
END OAI22X2H7R

MACRO OAI22X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22X3H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 2.025 1.095 2.165 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 0.795 -0.08 0.935 0.335 ;
        RECT 0.295 -0.08 0.435 0.335 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.195 0.655 0.535 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.695 0.655 1.035 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.885 0.655 2.225 0.745 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.505 0.655 1.775 0.765 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.325 0.425 2.125 0.515 ;
        RECT 1.985 0.35 2.125 0.515 ;
        RECT 1.525 0.855 1.665 1.02 ;
        RECT 0.795 0.855 1.665 0.945 ;
        RECT 1.325 0.35 1.465 0.515 ;
        RECT 1.325 0.35 1.415 0.945 ;
        RECT 0.795 0.855 0.935 1.02 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.275 1.11 1.89 1.2 ;
      RECT 1.8 0.915 1.89 1.2 ;
      RECT 1.275 1.08 1.415 1.2 ;
      RECT 2.275 0.915 2.415 1.035 ;
      RECT 1.8 0.915 2.415 1.005 ;
      RECT 0.07 0.425 1.16 0.515 ;
      RECT 1.07 0.17 1.16 0.515 ;
      RECT 0.57 0.295 0.66 0.515 ;
      RECT 0.07 0.28 0.16 0.515 ;
      RECT 2.29 0.17 2.38 0.395 ;
      RECT 1.605 0.17 1.745 0.335 ;
      RECT 1.07 0.17 2.38 0.26 ;
      RECT 0.57 1.11 1.185 1.2 ;
      RECT 1.045 1.08 1.185 1.2 ;
      RECT 0.57 0.905 0.66 1.2 ;
      RECT 0.07 0.905 0.16 1.06 ;
      RECT 0.07 0.905 0.66 0.995 ;
  END
END OAI22X3H7R

MACRO OAI22X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22X4H7R 0 0 ;
  SIZE 3 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3 1.48 ;
        RECT 2.277 1.095 2.417 1.48 ;
        RECT 0.547 1.095 0.687 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3 0.08 ;
        RECT 1.047 -0.08 1.187 0.305 ;
        RECT 0.547 -0.08 0.687 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.477 0.655 0.817 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.977 0.655 1.317 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.137 0.655 2.477 0.745 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.802 0.595 1.952 0.775 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.577 0.395 2.347 0.485 ;
        RECT 1.047 0.885 1.917 0.975 ;
        RECT 1.047 0.855 1.667 0.975 ;
        RECT 1.577 0.395 1.667 0.975 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.527 1.065 2.142 1.155 ;
      RECT 2.052 0.915 2.142 1.155 ;
      RECT 2.052 0.915 2.667 1.005 ;
      RECT 0.322 0.395 1.367 0.485 ;
      RECT 1.277 0.215 1.367 0.485 ;
      RECT 0.322 0.345 0.412 0.485 ;
      RECT 2.482 0.215 2.572 0.355 ;
      RECT 1.277 0.215 2.572 0.305 ;
      RECT 0.822 1.065 1.437 1.155 ;
      RECT 0.822 0.905 0.912 1.155 ;
      RECT 0.297 0.905 0.912 0.995 ;
  END
END OAI22X4H7R

MACRO OAI22X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22X6H7R 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.8 1.48 ;
        RECT 3.322 0.855 3.412 1.48 ;
        RECT 2.822 1.07 2.912 1.48 ;
        RECT 0.797 1.095 0.937 1.48 ;
        RECT 0.322 0.855 0.412 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.8 0.08 ;
        RECT 1.547 -0.08 1.687 0.305 ;
        RECT 1.047 -0.08 1.187 0.305 ;
        RECT 0.547 -0.08 0.687 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.477 0.655 1.017 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.227 0.655 1.767 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.727 0.655 3.267 0.745 ;
      LAYER MET2 ;
        RECT 2.85 0.43 2.95 0.96 ;
      LAYER VIA1 ;
        RECT 2.855 0.655 2.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.365 0.625 2.59 0.745 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.047 0.395 3.187 0.485 ;
        RECT 1.297 0.885 2.437 0.975 ;
        RECT 2.055 0.395 2.145 0.975 ;
      LAYER MET2 ;
        RECT 2.05 0.63 2.15 1.16 ;
      LAYER VIA1 ;
        RECT 2.055 0.855 2.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.322 0.395 1.912 0.485 ;
      RECT 1.822 0.215 1.912 0.485 ;
      RECT 0.322 0.345 0.412 0.485 ;
      RECT 3.322 0.215 3.412 0.355 ;
      RECT 1.822 0.215 3.412 0.305 ;
      RECT 3.072 0.855 3.162 1.2 ;
      RECT 2.047 1.065 2.662 1.155 ;
      RECT 2.572 0.855 2.662 1.155 ;
      RECT 2.572 0.855 3.162 0.945 ;
      RECT 1.072 1.065 1.687 1.155 ;
      RECT 1.072 0.905 1.162 1.155 ;
      RECT 0.547 0.905 1.162 0.995 ;
  END
END OAI22X6H7R

MACRO OAI2BB1X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB1X0P5H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.13 1.2 1.22 1.48 ;
        RECT 0.6 1.2 0.69 1.48 ;
        RECT 0.07 1.2 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.575 -0.08 0.715 0.175 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.455 0.575 0.545 ;
        RECT 0.47 0.455 0.56 0.695 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.24 0.625 0.345 0.775 ;
        RECT 0.24 0.5 0.33 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.625 0.79 0.775 ;
        RECT 0.7 0.55 0.79 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.84 0.855 1.215 0.945 ;
        RECT 1.125 0.23 1.215 0.945 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.06 0.865 0.45 0.955 ;
      RECT 0.06 0.275 0.15 0.955 ;
      RECT 0.945 0.275 1.035 0.73 ;
      RECT 0.06 0.275 1.035 0.365 ;
  END
END OAI2BB1X0P5H7R

MACRO OAI2BB1X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB1X0P7H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.24 1.055 1.33 1.48 ;
        RECT 0.73 1.07 0.82 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.715 -0.08 0.805 0.33 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.61 0.775 0.745 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.405 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.835 0.6 0.985 0.78 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.99 0.87 1.345 0.96 ;
        RECT 1.255 0.245 1.345 0.96 ;
        RECT 1.2 0.245 1.345 0.335 ;
        RECT 0.99 0.87 1.08 1.108 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.375 0.865 0.465 1.14 ;
      RECT 0.045 0.865 0.465 0.955 ;
      RECT 0.045 0.23 0.135 0.955 ;
      RECT 1.075 0.42 1.165 0.58 ;
      RECT 0.485 0.42 1.165 0.51 ;
      RECT 0.485 0.23 0.575 0.51 ;
      RECT 0.045 0.23 0.575 0.32 ;
  END
END OAI2BB1X0P7H7R

MACRO OAI2BB1X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB1X1H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.13 1.2 1.22 1.48 ;
        RECT 0.6 1.2 0.69 1.48 ;
        RECT 0.07 1.2 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.575 -0.08 0.715 0.175 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.455 0.575 0.545 ;
        RECT 0.465 0.455 0.555 0.695 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.655 0.375 0.745 ;
        RECT 0.225 0.505 0.315 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.625 0.795 0.775 ;
        RECT 0.675 0.575 0.795 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.84 0.855 1.215 0.945 ;
        RECT 1.125 0.285 1.215 0.945 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.835 0.45 0.925 ;
      RECT 0.045 0.265 0.135 0.925 ;
      RECT 0.945 0.265 1.035 0.695 ;
      RECT 0.045 0.265 1.035 0.355 ;
  END
END OAI2BB1X1H7R

MACRO OAI2BB1X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB1X1P4H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.215 1.08 1.355 1.48 ;
        RECT 0.73 1.07 0.82 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.715 -0.08 0.805 0.33 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.615 0.825 0.745 0.975 ;
        RECT 0.615 0.68 0.705 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.595 0.375 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.835 0.62 0.985 0.8 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.99 0.9 1.345 0.99 ;
        RECT 1.255 0.26 1.345 0.99 ;
        RECT 1.2 0.26 1.345 0.35 ;
        RECT 0.99 0.9 1.08 1.04 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.375 0.865 0.465 1.14 ;
      RECT 0.045 0.865 0.465 0.955 ;
      RECT 0.045 0.23 0.135 0.955 ;
      RECT 1.075 0.44 1.165 0.65 ;
      RECT 0.485 0.44 1.165 0.53 ;
      RECT 0.485 0.23 0.575 0.53 ;
      RECT 0.045 0.23 0.575 0.32 ;
  END
END OAI2BB1X1P4H7R

MACRO OAI2BB1X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB1X2H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.145 1.055 1.235 1.48 ;
        RECT 0.635 1.07 0.725 1.48 ;
        RECT 0.045 1.19 0.185 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.565 -0.08 0.655 0.33 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.435 0.75 0.555 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.615 0.345 0.84 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.615 0.805 0.795 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.895 0.855 1.265 0.945 ;
        RECT 1.175 0.255 1.265 0.945 ;
        RECT 1.07 0.255 1.265 0.345 ;
        RECT 0.895 0.855 0.985 1.195 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.281 1.065 0.5 1.155 ;
      RECT 0.273 1.023 0.281 1.151 ;
      RECT 0.227 0.996 0.273 1.124 ;
      RECT 0.181 0.95 0.227 1.078 ;
      RECT 0.181 1.046 0.319 1.078 ;
      RECT 0.135 0.904 0.181 1.032 ;
      RECT 0.091 0.23 0.135 0.987 ;
      RECT 0.045 0.23 0.135 0.942 ;
      RECT 0.995 0.435 1.085 0.705 ;
      RECT 0.36 0.435 1.085 0.525 ;
      RECT 0.36 0.23 0.45 0.525 ;
      RECT 0.045 0.23 0.45 0.32 ;
  END
END OAI2BB1X2H7R

MACRO OAI2BB1X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB1X3H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.63 1.08 1.77 1.48 ;
        RECT 1.145 1.07 1.235 1.48 ;
        RECT 0.635 1.07 0.725 1.48 ;
        RECT 0.045 1.195 0.185 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.055 -0.08 1.195 0.19 ;
        RECT 0.565 -0.08 0.655 0.35 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.705 0.555 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.36 0.825 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.72 0.655 1.06 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.895 0.855 1.82 0.945 ;
        RECT 1.73 0.449 1.82 0.945 ;
        RECT 1.631 0.404 1.776 0.463 ;
        RECT 1.55 0.365 1.73 0.44 ;
        RECT 1.699 0.449 1.82 0.524 ;
        RECT 1.55 0.35 1.699 0.44 ;
        RECT 1.677 0.449 1.82 0.497 ;
        RECT 1.405 0.855 1.495 1.045 ;
        RECT 0.895 0.855 0.985 1.045 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.79 0.28 1.4 0.37 ;
      RECT 1.31 0.17 1.4 0.37 ;
      RECT 1.84 0.17 1.93 0.345 ;
      RECT 1.31 0.17 1.93 0.26 ;
      RECT 0.276 1.065 0.5 1.155 ;
      RECT 0.273 1.025 0.276 1.154 ;
      RECT 0.227 1.001 0.273 1.129 ;
      RECT 0.181 0.955 0.227 1.083 ;
      RECT 0.181 1.046 0.314 1.083 ;
      RECT 0.135 0.909 0.181 1.037 ;
      RECT 0.091 0.31 0.135 0.992 ;
      RECT 0.045 0.31 0.135 0.947 ;
      RECT 1.3 0.64 1.64 0.73 ;
      RECT 1.3 0.46 1.39 0.73 ;
      RECT 0.476 0.46 1.39 0.55 ;
      RECT 0.456 0.412 0.476 0.54 ;
      RECT 0.41 0.379 0.456 0.507 ;
      RECT 0.364 0.333 0.41 0.461 ;
      RECT 0.364 0.441 0.514 0.461 ;
      RECT 0.326 0.31 0.364 0.419 ;
      RECT 0.045 0.31 0.364 0.4 ;
  END
END OAI2BB1X3H7R

MACRO OAI2BB1X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB1X4H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 1.655 1.055 1.745 1.48 ;
        RECT 1.145 1.07 1.235 1.48 ;
        RECT 0.635 1.07 0.725 1.48 ;
        RECT 0.045 1.19 0.185 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 1.105 -0.08 1.245 0.175 ;
        RECT 0.565 -0.08 0.655 0.33 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.685 0.555 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.36 0.825 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.72 0.655 1.06 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.895 0.855 1.82 0.945 ;
        RECT 1.73 0.418 1.82 0.945 ;
        RECT 1.585 0.395 1.774 0.485 ;
        RECT 0.895 0.855 0.985 1 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END Z
  OBS
    LAYER MET1 ;
      RECT 0.79 0.265 1.45 0.355 ;
      RECT 1.36 0.17 1.45 0.355 ;
      RECT 1.86 0.17 1.95 0.345 ;
      RECT 1.36 0.17 1.95 0.26 ;
      RECT 0.281 1.065 0.5 1.155 ;
      RECT 0.273 1.023 0.281 1.151 ;
      RECT 0.227 0.996 0.273 1.124 ;
      RECT 0.181 0.95 0.227 1.078 ;
      RECT 0.181 1.046 0.319 1.078 ;
      RECT 0.135 0.904 0.181 1.032 ;
      RECT 0.091 0.25 0.135 0.987 ;
      RECT 0.045 0.25 0.135 0.942 ;
      RECT 1.3 0.625 1.64 0.715 ;
      RECT 1.3 0.445 1.39 0.715 ;
      RECT 0.36 0.445 1.39 0.535 ;
      RECT 0.36 0.25 0.45 0.535 ;
      RECT 0.045 0.25 0.45 0.34 ;
  END
END OAI2BB1X4H7R

MACRO OAI2BB1X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB1X6H7R 0 0 ;
  SIZE 2.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.8 1.48 ;
        RECT 2.345 1.08 2.485 1.48 ;
        RECT 1.87 1.07 1.96 1.48 ;
        RECT 1.36 1.07 1.45 1.48 ;
        RECT 0.85 1.07 0.94 1.48 ;
        RECT 0.26 1.19 0.4 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.8 0.08 ;
        RECT 1.32 -0.08 1.46 0.175 ;
        RECT 0.78 -0.08 0.87 0.33 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.615 0.77 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.615 0.56 0.84 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.935 0.655 1.475 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.885 0.395 2.5 0.485 ;
        RECT 2.41 0.315 2.5 0.485 ;
        RECT 1.085 0.885 2.345 0.975 ;
        RECT 2.255 0.395 2.345 0.975 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.005 0.265 1.75 0.355 ;
      RECT 1.66 0.17 1.75 0.355 ;
      RECT 2.135 0.17 2.275 0.305 ;
      RECT 1.66 0.17 2.275 0.26 ;
      RECT 0.496 1.065 0.715 1.155 ;
      RECT 0.488 1.023 0.496 1.151 ;
      RECT 0.442 0.996 0.488 1.124 ;
      RECT 0.396 0.95 0.442 1.078 ;
      RECT 0.396 1.046 0.534 1.078 ;
      RECT 0.35 0.904 0.396 1.032 ;
      RECT 0.306 0.345 0.35 0.987 ;
      RECT 0.26 0.345 0.35 0.942 ;
      RECT 1.705 0.655 2.115 0.745 ;
      RECT 1.705 0.445 1.795 0.745 ;
      RECT 0.835 0.445 1.795 0.535 ;
      RECT 0.575 0.435 0.925 0.525 ;
      RECT 0.26 0.345 0.665 0.435 ;
  END
END OAI2BB1X6H7R

MACRO OAI2BB2X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB2X0P5H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.335 1.24 1.475 1.48 ;
        RECT 0.57 1.07 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.03 -0.08 1.17 0.32 ;
        RECT 0.555 -0.08 0.645 0.33 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.55 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.425 0.545 0.695 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.595 0.805 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.905 0.645 1.175 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.005 1.055 1.625 1.145 ;
        RECT 1.535 0.205 1.625 1.145 ;
      LAYER MET2 ;
        RECT 1.45 0.84 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.805 0.41 1.375 0.5 ;
      RECT 1.285 0.205 1.375 0.5 ;
      RECT 0.805 0.22 0.895 0.5 ;
      RECT 0.32 0.865 0.41 1.14 ;
      RECT 0.045 0.865 1.325 0.955 ;
      RECT 1.235 0.815 1.325 0.955 ;
      RECT 0.045 0.23 0.135 0.955 ;
      RECT 0.045 0.23 0.185 0.32 ;
  END
END OAI2BB2X0P5H7R

MACRO OAI2BB2X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB2X0P7H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.335 1.235 1.475 1.48 ;
        RECT 0.57 1.07 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.03 -0.08 1.17 0.32 ;
        RECT 0.555 -0.08 0.645 0.33 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.545 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.435 0.425 0.555 0.65 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.595 0.805 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.905 0.645 1.175 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.005 1.055 1.625 1.145 ;
        RECT 1.535 0.23 1.625 1.145 ;
      LAYER MET2 ;
        RECT 1.45 0.84 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.805 0.41 1.375 0.5 ;
      RECT 1.285 0.23 1.375 0.5 ;
      RECT 0.805 0.245 0.895 0.5 ;
      RECT 0.32 0.865 0.41 1.14 ;
      RECT 0.045 0.865 1.34 0.955 ;
      RECT 1.25 0.795 1.34 0.955 ;
      RECT 0.045 0.23 0.135 0.955 ;
      RECT 0.045 0.23 0.185 0.32 ;
  END
END OAI2BB2X0P7H7R

MACRO OAI2BB2X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB2X1H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.335 1.235 1.475 1.48 ;
        RECT 0.57 1.07 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.03 -0.08 1.17 0.32 ;
        RECT 0.555 -0.08 0.645 0.33 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.55 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.435 0.425 0.555 0.65 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.595 0.805 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.905 0.645 1.175 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.005 1.055 1.625 1.145 ;
        RECT 1.535 0.265 1.625 1.145 ;
      LAYER MET2 ;
        RECT 1.45 0.84 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.805 0.41 1.375 0.5 ;
      RECT 1.285 0.265 1.375 0.5 ;
      RECT 0.805 0.28 0.895 0.5 ;
      RECT 0.32 0.865 0.41 1.14 ;
      RECT 0.045 0.865 1.355 0.955 ;
      RECT 1.265 0.75 1.355 0.955 ;
      RECT 0.045 0.23 0.135 0.955 ;
      RECT 0.045 0.23 0.185 0.32 ;
  END
END OAI2BB2X1H7R

MACRO OAI2BB2X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB2X1P4H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.335 1.235 1.475 1.48 ;
        RECT 0.57 1.07 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.03 -0.08 1.17 0.32 ;
        RECT 0.555 -0.08 0.645 0.33 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.55 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.435 0.425 0.555 0.65 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.595 0.805 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.905 0.645 1.175 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.005 1.055 1.625 1.145 ;
        RECT 1.535 0.3 1.625 1.145 ;
      LAYER MET2 ;
        RECT 1.45 0.84 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.805 0.41 1.375 0.5 ;
      RECT 1.285 0.3 1.375 0.5 ;
      RECT 0.805 0.315 0.895 0.5 ;
      RECT 0.32 0.865 0.41 1.14 ;
      RECT 0.045 0.865 1.355 0.955 ;
      RECT 1.265 0.705 1.355 0.955 ;
      RECT 0.045 0.23 0.135 0.955 ;
      RECT 0.045 0.23 0.185 0.32 ;
  END
END OAI2BB2X1P4H7R

MACRO OAI2BB2X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB2X2H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.335 1.235 1.475 1.48 ;
        RECT 0.57 1.07 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.03 -0.08 1.17 0.32 ;
        RECT 0.555 -0.08 0.645 0.33 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.55 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.425 0.545 0.725 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.595 0.805 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.915 0.64 1.175 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.005 1.055 1.625 1.145 ;
        RECT 1.535 0.355 1.625 1.145 ;
      LAYER MET2 ;
        RECT 1.45 0.84 1.55 1.22 ;
      LAYER VIA1 ;
        RECT 1.455 1.055 1.545 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.805 0.41 1.375 0.5 ;
      RECT 1.285 0.355 1.375 0.5 ;
      RECT 0.805 0.36 0.895 0.5 ;
      RECT 0.32 0.865 0.41 1.14 ;
      RECT 0.045 0.865 1.355 0.955 ;
      RECT 1.265 0.64 1.355 0.955 ;
      RECT 0.045 0.23 0.135 0.955 ;
      RECT 0.045 0.23 0.185 0.32 ;
  END
END OAI2BB2X2H7R

MACRO OAI2BB2X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB2X3H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 2.155 1.095 2.295 1.48 ;
        RECT 1.11 1.225 1.25 1.48 ;
        RECT 0.57 1.07 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 1.595 -0.08 1.735 0.175 ;
        RECT 1.03 -0.08 1.17 0.305 ;
        RECT 0.555 -0.08 0.645 0.33 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.55 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.425 0.545 0.725 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.68 0.655 1.02 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.485 0.49 1.825 0.58 ;
        RECT 1.625 0.455 1.825 0.58 ;
      LAYER MET2 ;
        RECT 1.65 0.23 1.75 0.76 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.43 0.915 2.545 1.06 ;
        RECT 2.455 0.41 2.545 1.06 ;
        RECT 2.1 0.41 2.545 0.5 ;
        RECT 1.93 0.915 2.545 1.005 ;
        RECT 2.1 0.35 2.24 0.5 ;
        RECT 1.34 1.11 2.02 1.2 ;
        RECT 1.93 0.915 2.02 1.2 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.805 0.395 1.395 0.485 ;
      RECT 1.305 0.265 1.395 0.485 ;
      RECT 0.805 0.295 0.895 0.485 ;
      RECT 1.305 0.265 1.94 0.355 ;
      RECT 1.85 0.17 1.94 0.355 ;
      RECT 2.365 0.17 2.505 0.32 ;
      RECT 1.85 0.17 2.505 0.26 ;
      RECT 0.32 0.865 0.41 1.06 ;
      RECT 0.045 0.865 1.102 0.955 ;
      RECT 0.045 0.865 1.148 0.932 ;
      RECT 1.064 0.846 1.194 0.886 ;
      RECT 0.045 0.29 0.135 0.955 ;
      RECT 1.102 0.804 1.194 0.886 ;
      RECT 1.102 0.804 1.232 0.844 ;
      RECT 1.194 0.735 2.355 0.825 ;
      RECT 1.148 0.758 2.355 0.825 ;
      RECT 0.045 0.29 0.185 0.38 ;
      RECT 0.795 1.045 1.178 1.135 ;
      RECT 0.795 1.045 1.224 1.112 ;
      RECT 1.14 1.026 1.255 1.074 ;
      RECT 1.178 0.984 1.293 1.039 ;
      RECT 1.224 0.945 1.255 1.074 ;
      RECT 1.255 0.93 1.795 1.02 ;
  END
END OAI2BB2X3H7R

MACRO OAI2BB2X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB2X4H7R 0 0 ;
  SIZE 2.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.8 1.48 ;
        RECT 2.155 1.095 2.295 1.48 ;
        RECT 1.11 1.225 1.25 1.48 ;
        RECT 0.57 1.07 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.8 0.08 ;
        RECT 1.595 -0.08 1.735 0.175 ;
        RECT 1.03 -0.08 1.17 0.305 ;
        RECT 0.555 -0.08 0.645 0.33 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.55 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.425 0.545 0.725 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.71 0.655 1.05 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.459 0.565 1.799 0.655 ;
        RECT 1.625 0.455 1.799 0.655 ;
      LAYER MET2 ;
        RECT 1.65 0.23 1.75 0.76 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.93 0.915 2.545 1.005 ;
        RECT 2.455 0.41 2.545 1.005 ;
        RECT 2.085 0.41 2.545 0.5 ;
        RECT 2.085 0.395 2.225 0.5 ;
        RECT 1.34 1.105 2.02 1.195 ;
        RECT 1.93 0.915 2.02 1.195 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.78 0.395 1.395 0.485 ;
      RECT 1.305 0.265 1.395 0.485 ;
      RECT 1.305 0.265 1.94 0.355 ;
      RECT 2.335 0.215 2.475 0.32 ;
      RECT 1.85 0.215 2.475 0.305 ;
      RECT 0.32 0.865 0.41 1.02 ;
      RECT 0.045 0.865 1.102 0.955 ;
      RECT 0.045 0.865 1.148 0.932 ;
      RECT 1.064 0.846 1.184 0.891 ;
      RECT 0.045 0.33 0.135 0.955 ;
      RECT 1.102 0.804 1.222 0.854 ;
      RECT 1.102 0.804 1.886 0.835 ;
      RECT 1.148 0.763 1.928 0.814 ;
      RECT 1.184 0.745 1.966 0.774 ;
      RECT 1.886 0.686 1.928 0.814 ;
      RECT 1.928 0.665 2.355 0.755 ;
      RECT 1.848 0.726 2.355 0.755 ;
      RECT 0.045 0.33 0.185 0.42 ;
      RECT 0.795 1.045 1.178 1.135 ;
      RECT 0.795 1.045 1.224 1.112 ;
      RECT 1.14 1.026 1.26 1.071 ;
      RECT 1.178 0.984 1.298 1.034 ;
      RECT 1.224 0.943 1.26 1.071 ;
      RECT 1.26 0.925 1.795 1.015 ;
  END
END OAI2BB2X4H7R

MACRO OAI2BB2X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB2X6H7R 0 0 ;
  SIZE 4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4 1.48 ;
        RECT 3.295 0.855 3.385 1.48 ;
        RECT 2.795 1.07 2.885 1.48 ;
        RECT 1.325 1.225 1.465 1.48 ;
        RECT 0.785 1.07 0.875 1.48 ;
        RECT 0.285 1.055 0.375 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4 0.08 ;
        RECT 2.385 -0.08 2.525 0.185 ;
        RECT 1.82 -0.08 1.96 0.305 ;
        RECT 1.245 -0.08 1.385 0.305 ;
        RECT 0.745 -0.08 0.885 0.305 ;
    END
  END VSS
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.55 0.56 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.425 0.76 0.705 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.925 0.655 1.265 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.14 0.565 2.48 0.655 ;
        RECT 2.225 0.455 2.375 0.655 ;
      LAYER MET2 ;
        RECT 2.25 0.23 2.35 0.76 ;
      LAYER VIA1 ;
        RECT 2.255 0.455 2.345 0.545 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.875 0.395 3.49 0.485 ;
        RECT 3.4 0.345 3.49 0.485 ;
        RECT 3.115 0.395 3.205 0.945 ;
        RECT 2.681 0.892 3.205 0.945 ;
        RECT 2.741 0.855 3.205 0.945 ;
        RECT 2.635 0.938 2.779 0.964 ;
        RECT 2.635 0.938 2.741 0.99 ;
        RECT 2.727 0.862 3.205 0.945 ;
        RECT 2.591 0.983 2.727 1.02 ;
        RECT 2.591 0.983 2.681 1.066 ;
        RECT 1.955 1.105 2.635 1.195 ;
        RECT 2.545 1.028 2.635 1.195 ;
      LAYER MET2 ;
        RECT 3.05 0.63 3.15 1.16 ;
      LAYER VIA1 ;
        RECT 3.055 0.855 3.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.995 0.395 2.039 0.485 ;
      RECT 2.001 0.376 2.116 0.431 ;
      RECT 2.039 0.341 2.07 0.47 ;
      RECT 2.07 0.275 2.159 0.387 ;
      RECT 2.07 0.275 2.73 0.365 ;
      RECT 2.64 0.215 3.265 0.305 ;
      RECT 0.26 0.865 1.575 0.955 ;
      RECT 1.485 0.745 1.575 0.955 ;
      RECT 0.26 0.355 0.35 0.955 ;
      RECT 1.485 0.745 2.631 0.835 ;
      RECT 1.485 0.745 2.677 0.812 ;
      RECT 1.485 0.745 2.721 0.764 ;
      RECT 2.683 0.655 3.025 0.745 ;
      RECT 2.593 0.726 3.025 0.745 ;
      RECT 2.677 0.658 2.683 0.786 ;
      RECT 2.631 0.684 3.025 0.745 ;
      RECT 0.26 0.355 0.4 0.445 ;
      RECT 1.01 1.045 1.755 1.135 ;
      RECT 1.665 0.925 1.755 1.135 ;
      RECT 1.665 0.925 2.41 1.015 ;
  END
END OAI2BB2X6H7R

MACRO OAI2XB1X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2XB1X0P5H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.985 1.095 1.125 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.775 -0.08 0.915 0.305 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.605 1.005 0.785 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A0
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.165 0.625 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.165 0.625 1.345 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.74 0.915 1.545 1.005 ;
        RECT 1.455 0.23 1.545 1.005 ;
        RECT 1.275 0.23 1.545 0.32 ;
        RECT 1.26 0.915 1.35 1.155 ;
        RECT 0.525 1.045 0.83 1.135 ;
        RECT 0.74 0.915 0.83 1.135 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.686 0.395 1.14 0.485 ;
      RECT 1.05 0.22 1.14 0.485 ;
      RECT 0.64 0.334 0.686 0.462 ;
      RECT 0.596 0.205 0.64 0.417 ;
      RECT 0.596 0.376 0.724 0.417 ;
      RECT 0.55 0.205 0.64 0.372 ;
      RECT 0.32 0.865 0.41 1.155 ;
      RECT 0.32 0.865 0.525 0.955 ;
      RECT 0.435 0.509 0.525 0.955 ;
      RECT 0.435 0.635 0.735 0.725 ;
      RECT 0.41 0.428 0.435 0.557 ;
      RECT 0.366 0.464 0.481 0.522 ;
      RECT 0.32 0.205 0.41 0.477 ;
  END
END OAI2XB1X0P5H7R

MACRO OAI2XB1X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2XB1X0P7H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.985 1.095 1.125 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.775 -0.08 0.915 0.305 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.605 1.005 0.785 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A0
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.165 0.625 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.165 0.625 1.345 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.645 0.915 1.545 1.005 ;
        RECT 1.455 0.254 1.545 1.005 ;
        RECT 1.275 0.254 1.545 0.344 ;
        RECT 1.26 0.915 1.35 1.125 ;
        RECT 0.525 1.045 0.735 1.135 ;
        RECT 0.645 0.915 0.735 1.135 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.646 0.395 1.14 0.485 ;
      RECT 1.05 0.244 1.14 0.485 ;
      RECT 0.64 0.354 0.646 0.482 ;
      RECT 0.596 0.395 1.14 0.457 ;
      RECT 0.55 0.229 0.64 0.412 ;
      RECT 0.55 0.376 0.684 0.412 ;
      RECT 0.32 0.865 0.41 1.155 ;
      RECT 0.32 0.865 0.525 0.955 ;
      RECT 0.435 0.489 0.525 0.955 ;
      RECT 0.435 0.635 0.735 0.725 ;
      RECT 0.41 0.408 0.435 0.537 ;
      RECT 0.366 0.444 0.481 0.502 ;
      RECT 0.32 0.205 0.41 0.457 ;
  END
END OAI2XB1X0P7H7R

MACRO OAI2XB1X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2XB1X1H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.985 1.095 1.125 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.775 -0.08 0.915 0.305 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.605 1.005 0.785 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A0
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.165 0.625 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.165 0.625 1.345 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.915 1.545 1.005 ;
        RECT 1.455 0.29 1.545 1.005 ;
        RECT 1.275 0.29 1.545 0.38 ;
        RECT 1.26 0.915 1.35 1.075 ;
        RECT 0.525 1.045 0.745 1.135 ;
        RECT 0.655 0.915 0.745 1.135 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.626 0.395 1.14 0.485 ;
      RECT 1.05 0.28 1.14 0.485 ;
      RECT 0.596 0.395 1.14 0.47 ;
      RECT 0.55 0.265 0.64 0.432 ;
      RECT 0.55 0.383 0.664 0.432 ;
      RECT 0.32 0.865 0.41 1.155 ;
      RECT 0.32 0.865 0.525 0.955 ;
      RECT 0.435 0.504 0.525 0.955 ;
      RECT 0.435 0.635 0.735 0.725 ;
      RECT 0.41 0.423 0.435 0.552 ;
      RECT 0.366 0.459 0.481 0.517 ;
      RECT 0.32 0.205 0.41 0.472 ;
  END
END OAI2XB1X1H7R

MACRO OAI2XB1X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2XB1X1P4H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.985 1.095 1.125 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.775 -0.08 0.915 0.305 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.6 1.005 0.78 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A0
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.165 0.625 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.11 0.58 1.345 0.79 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.915 1.545 1.005 ;
        RECT 1.455 0.326 1.545 1.005 ;
        RECT 1.275 0.326 1.545 0.416 ;
        RECT 0.525 1.045 0.745 1.135 ;
        RECT 0.655 0.915 0.745 1.135 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.596 0.395 1.14 0.485 ;
      RECT 1.05 0.316 1.14 0.485 ;
      RECT 0.55 0.295 0.64 0.462 ;
      RECT 0.32 0.865 0.41 1.155 ;
      RECT 0.32 0.865 0.525 0.955 ;
      RECT 0.435 0.524 0.525 0.955 ;
      RECT 0.435 0.635 0.735 0.725 ;
      RECT 0.41 0.443 0.435 0.572 ;
      RECT 0.366 0.479 0.481 0.537 ;
      RECT 0.32 0.205 0.41 0.492 ;
  END
END OAI2XB1X1P4H7R

MACRO OAI2XB1X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2XB1X2H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.01 1.07 1.1 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 0.775 -0.08 0.915 0.305 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.605 1.005 0.785 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A0
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.165 0.625 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.17 0.615 1.345 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.65 0.885 1.545 0.975 ;
        RECT 1.455 0.38 1.545 0.975 ;
        RECT 1.275 0.38 1.545 0.47 ;
        RECT 0.525 1.045 0.74 1.135 ;
        RECT 0.65 0.885 0.74 1.135 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.596 0.395 1.165 0.485 ;
      RECT 0.55 0.295 0.64 0.462 ;
      RECT 0.32 0.865 0.41 1.155 ;
      RECT 0.32 0.865 0.525 0.955 ;
      RECT 0.435 0.524 0.525 0.955 ;
      RECT 0.435 0.635 0.735 0.725 ;
      RECT 0.41 0.443 0.435 0.572 ;
      RECT 0.366 0.479 0.481 0.537 ;
      RECT 0.32 0.205 0.41 0.492 ;
  END
END OAI2XB1X2H7R

MACRO OAI2XB1X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2XB1X3H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 2.345 1.055 2.435 1.48 ;
        RECT 1.845 1.07 1.935 1.48 ;
        RECT 1.255 1.215 1.395 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 1.5 -0.08 1.64 0.305 ;
        RECT 0.775 -0.08 0.915 0.305 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.24 0.655 1.78 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A0
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.165 0.625 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.165 0.625 2.345 0.775 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.053 0.93 2.21 1.02 ;
        RECT 1.985 0.35 2.17 0.44 ;
        RECT 0.879 0.922 2.091 0.945 ;
        RECT 0.879 0.911 2.075 0.945 ;
        RECT 2.031 0.93 2.21 1.009 ;
        RECT 1.985 0.35 2.075 0.975 ;
        RECT 1.978 0.93 2.21 0.949 ;
        RECT 0.917 0.873 2.075 0.945 ;
        RECT 0.954 0.855 2.075 0.945 ;
        RECT 0.775 0.93 0.992 0.964 ;
        RECT 0.775 0.93 0.954 1.002 ;
        RECT 0.775 0.93 0.917 1.02 ;
      LAYER MET2 ;
        RECT 1.85 0.625 1.95 1.16 ;
      LAYER VIA1 ;
        RECT 1.855 0.855 1.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.615 0.395 1.865 0.485 ;
      RECT 1.775 0.17 1.865 0.485 ;
      RECT 0.596 0.395 1.865 0.476 ;
      RECT 0.55 0.28 0.64 0.443 ;
      RECT 1.155 0.295 1.245 0.485 ;
      RECT 0.55 0.388 0.653 0.443 ;
      RECT 2.335 0.17 2.425 0.345 ;
      RECT 1.775 0.17 2.425 0.26 ;
      RECT 0.55 1.11 1.14 1.2 ;
      RECT 1.05 1.035 1.71 1.125 ;
      RECT 0.55 1.055 0.64 1.2 ;
      RECT 0.32 0.865 0.41 1.155 ;
      RECT 0.32 0.865 0.57 0.955 ;
      RECT 0.48 0.575 0.57 0.955 ;
      RECT 0.48 0.575 0.985 0.665 ;
      RECT 0.456 0.474 0.48 0.602 ;
      RECT 0.456 0.553 0.569 0.602 ;
      RECT 0.41 0.439 0.456 0.567 ;
      RECT 0.41 0.509 0.526 0.567 ;
      RECT 0.366 0.265 0.41 0.522 ;
      RECT 0.32 0.265 0.41 0.477 ;
  END
END OAI2XB1X3H7R

MACRO OAI2XB1X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2XB1X4H7R 0 0 ;
  SIZE 2.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.8 1.48 ;
        RECT 2.345 1.055 2.435 1.48 ;
        RECT 1.845 1.07 1.935 1.48 ;
        RECT 1.255 1.215 1.395 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.8 0.08 ;
        RECT 1.5 -0.08 1.64 0.305 ;
        RECT 0.775 -0.08 0.915 0.305 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.24 0.655 1.78 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A0
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.165 0.625 0.345 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.165 0.625 2.345 0.775 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.985 0.885 2.21 0.975 ;
        RECT 1.985 0.35 2.14 0.44 ;
        RECT 0.775 0.855 2.075 0.945 ;
        RECT 1.985 0.35 2.075 0.975 ;
      LAYER MET2 ;
        RECT 1.85 0.625 1.95 1.16 ;
      LAYER VIA1 ;
        RECT 1.855 0.855 1.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.6 0.395 1.865 0.485 ;
      RECT 1.775 0.17 1.865 0.485 ;
      RECT 0.596 0.395 1.865 0.483 ;
      RECT 0.55 0.295 0.64 0.458 ;
      RECT 2.335 0.17 2.425 0.345 ;
      RECT 1.775 0.17 2.425 0.26 ;
      RECT 0.32 0.908 0.41 1.075 ;
      RECT 0.435 0.479 0.481 0.921 ;
      RECT 0.366 0.863 0.481 0.921 ;
      RECT 0.41 0.828 0.435 0.957 ;
      RECT 0.435 0.524 0.525 0.876 ;
      RECT 0.435 0.575 0.985 0.665 ;
      RECT 0.41 0.443 0.435 0.572 ;
      RECT 0.366 0.305 0.41 0.537 ;
      RECT 0.32 0.305 0.41 0.492 ;
      RECT 0.525 1.035 1.71 1.125 ;
  END
END OAI2XB1X4H7R

MACRO OAI2XB1X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2XB1X6H7R 0 0 ;
  SIZE 3.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.6 1.48 ;
        RECT 3.102 0.855 3.192 1.48 ;
        RECT 2.602 1.07 2.692 1.48 ;
        RECT 1.327 1.095 1.467 1.48 ;
        RECT 0.852 1.095 0.942 1.48 ;
        RECT 0.602 1.095 0.942 1.185 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.6 0.08 ;
        RECT 2.077 -0.08 2.217 0.305 ;
        RECT 1.577 -0.08 1.717 0.305 ;
        RECT 1.077 -0.08 1.217 0.305 ;
        RECT 0.555 -0.08 0.645 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.585 0.655 0.785 0.79 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A0
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.22 0.645 0.49 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.697 0.655 3.037 0.745 ;
      LAYER MET2 ;
        RECT 2.85 0.43 2.95 0.96 ;
      LAYER VIA1 ;
        RECT 2.855 0.655 2.945 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.487 0.395 3.217 0.485 ;
        RECT 3.077 0.38 3.217 0.485 ;
        RECT 1.827 0.885 2.967 0.975 ;
        RECT 1.827 0.855 2.577 0.975 ;
        RECT 2.487 0.395 2.577 0.975 ;
      LAYER MET2 ;
        RECT 2.45 0.625 2.55 1.16 ;
      LAYER VIA1 ;
        RECT 2.455 0.855 2.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.001 0.395 2.397 0.485 ;
      RECT 2.307 0.215 2.397 0.485 ;
      RECT 0.988 0.35 1.001 0.479 ;
      RECT 0.942 0.321 0.988 0.449 ;
      RECT 0.907 0.205 0.942 0.409 ;
      RECT 0.907 0.376 1.039 0.409 ;
      RECT 0.861 0.205 0.942 0.368 ;
      RECT 0.852 0.205 0.942 0.345 ;
      RECT 2.307 0.215 2.967 0.305 ;
      RECT 0.305 0.855 0.395 1.195 ;
      RECT 0.305 0.88 0.987 0.97 ;
      RECT 0.897 0.577 0.987 0.97 ;
      RECT 0.897 0.625 2.297 0.715 ;
      RECT 0.894 0.507 0.897 0.636 ;
      RECT 0.894 0.612 1.013 0.636 ;
      RECT 0.848 0.483 0.894 0.611 ;
      RECT 0.848 0.532 0.943 0.611 ;
      RECT 0.81 0.532 0.943 0.569 ;
      RECT 0.305 0.46 0.848 0.55 ;
      RECT 0.305 0.335 0.395 0.55 ;
      RECT 1.602 1.065 2.217 1.155 ;
      RECT 1.602 0.905 1.692 1.155 ;
      RECT 1.077 0.905 1.692 0.995 ;
  END
END OAI2XB1X6H7R

MACRO OAI31X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31X0P5H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.13 1.055 1.22 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.56 -0.08 0.7 0.255 ;
        RECT 0.07 -0.08 0.16 0.445 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.395 0.615 0.545 0.795 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.825 0.775 1.05 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.82 0.645 1.09 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.88 0.855 1.27 0.945 ;
        RECT 1.18 0.305 1.27 0.945 ;
        RECT 0.88 0.855 0.97 1.14 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.295 0.345 0.965 0.435 ;
  END
END OAI31X0P5H7R

MACRO OAI31X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31X0P7H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.12 1.055 1.21 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.56 -0.08 0.7 0.255 ;
        RECT 0.07 -0.08 0.16 0.42 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.575 0.545 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.63 0.823 0.78 1.003 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.645 1.095 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.87 0.855 1.275 0.945 ;
        RECT 1.185 0.33 1.275 0.945 ;
        RECT 1.075 0.33 1.275 0.42 ;
        RECT 0.87 0.855 0.96 1.108 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.295 0.345 0.965 0.435 ;
  END
END OAI31X0P7H7R

MACRO OAI31X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31X1H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.13 1.055 1.22 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.56 -0.08 0.7 0.255 ;
        RECT 0.07 -0.08 0.16 0.385 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.715 0.56 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.625 0.79 0.825 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.625 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.88 0.875 1.345 0.965 ;
        RECT 1.24 0.305 1.345 0.965 ;
        RECT 0.88 0.875 0.97 1.06 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.295 0.345 0.965 0.435 ;
  END
END OAI31X1H7R

MACRO OAI31X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31X1P4H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.13 1.055 1.22 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.6 -0.08 0.69 0.34 ;
        RECT 0.07 -0.08 0.16 0.355 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.395 0.625 0.545 0.92 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.706 0.81 0.796 ;
        RECT 0.655 0.706 0.745 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.98 0.455 1.175 0.545 ;
        RECT 0.98 0.455 1.07 0.67 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.585 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.88 0.855 1.355 0.945 ;
        RECT 1.265 0.25 1.355 0.945 ;
        RECT 1.135 0.25 1.355 0.34 ;
        RECT 0.88 0.855 0.97 1.02 ;
      LAYER MET2 ;
        RECT 1.05 0.815 1.15 1.22 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.38 0.43 0.89 0.52 ;
      RECT 0.8 0.25 0.89 0.52 ;
      RECT 0.38 0.25 0.47 0.52 ;
      RECT 0.8 0.25 0.995 0.34 ;
      RECT 0.295 0.25 0.47 0.34 ;
  END
END OAI31X1P4H7R

MACRO OAI31X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31X2H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.343 1.055 1.433 1.48 ;
        RECT 0.283 0.855 0.373 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 0.823 -0.08 0.963 0.26 ;
        RECT 0.283 -0.08 0.373 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.223 0.645 0.493 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.615 0.745 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.625 1.048 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.225 0.55 1.345 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.865 1.525 0.955 ;
        RECT 1.435 0.305 1.525 0.955 ;
        RECT 1.423 0.305 1.525 0.445 ;
        RECT 1.055 0.865 1.145 1.205 ;
      LAYER MET2 ;
        RECT 1.05 0.84 1.15 1.22 ;
      LAYER VIA1 ;
        RECT 1.055 1.055 1.145 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.508 0.36 1.278 0.45 ;
  END
END OAI31X2H7R

MACRO OAI31X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31X3H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 1.915 1.24 2.055 1.48 ;
        RECT 0.785 1.24 0.925 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 1.37 -0.08 1.51 0.175 ;
        RECT 0.84 -0.08 0.98 0.175 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.685 0.455 1.025 0.61 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.7 1.345 0.79 ;
        RECT 0.45 0.625 0.545 0.79 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.22 0.88 1.55 0.97 ;
        RECT 1.46 0.69 1.55 0.97 ;
        RECT 0.22 0.855 0.375 0.97 ;
        RECT 0.22 0.69 0.31 0.97 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.84 0.655 2.18 0.745 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.045 1.06 2.335 1.15 ;
        RECT 1.66 0.455 2.04 0.545 ;
        RECT 1.9 0.35 2.04 0.545 ;
        RECT 1.66 0.455 1.75 1.15 ;
      LAYER MET2 ;
        RECT 1.85 0.225 1.95 0.76 ;
      LAYER VIA1 ;
        RECT 1.855 0.455 1.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.19 0.17 2.28 0.375 ;
      RECT 0.045 0.275 1.75 0.365 ;
      RECT 1.66 0.17 1.75 0.365 ;
      RECT 1.66 0.17 2.28 0.26 ;
  END
END OAI31X3H7R

MACRO OAI31X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31X4H7R 0 0 ;
  SIZE 3.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.2 1.48 ;
        RECT 2.542 1.195 2.682 1.48 ;
        RECT 1.212 1.195 1.352 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.2 0.08 ;
        RECT 1.897 -0.08 2.037 0.175 ;
        RECT 1.267 -0.08 1.407 0.175 ;
        RECT 0.637 -0.08 0.777 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.175 0.655 1.515 0.745 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.707 0.455 1.797 0.705 ;
        RECT 0.797 0.455 1.797 0.545 ;
        RECT 0.797 0.455 0.887 0.68 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.835 2.162 0.925 ;
        RECT 2.072 0.615 2.162 0.925 ;
        RECT 0.455 0.615 0.599 0.925 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.432 0.655 2.808 0.745 ;
      LAYER MET2 ;
        RECT 2.65 0.43 2.75 0.96 ;
      LAYER VIA1 ;
        RECT 2.655 0.655 2.745 0.745 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.912 0.835 3.002 1.175 ;
        RECT 0.322 1.015 3.002 1.105 ;
        RECT 2.225 0.455 2.602 0.545 ;
        RECT 2.462 0.395 2.602 0.545 ;
        RECT 2.252 0.455 2.342 1.105 ;
      LAYER MET2 ;
        RECT 2.25 0.23 2.35 0.76 ;
      LAYER VIA1 ;
        RECT 2.255 0.455 2.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.322 0.275 2.327 0.365 ;
      RECT 2.737 0.215 2.827 0.355 ;
      RECT 2.237 0.215 2.827 0.305 ;
  END
END OAI31X4H7R

MACRO OAI32X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32X0P5H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.335 1.015 1.425 1.48 ;
        RECT 0.07 1.015 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.545 -0.08 0.685 0.36 ;
        RECT 0.07 -0.08 0.16 0.4 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.42 0.855 0.575 0.945 ;
        RECT 0.42 0.71 0.51 0.945 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.605 0.63 0.805 0.765 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.29 0.625 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.855 0.99 0.945 ;
        RECT 0.9 0.72 0.99 0.945 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.075 0.35 1.215 0.44 ;
        RECT 0.795 1.055 1.175 1.145 ;
        RECT 1.085 0.35 1.175 1.145 ;
      LAYER MET2 ;
        RECT 1.05 0.84 1.15 1.22 ;
      LAYER VIA1 ;
        RECT 1.055 1.055 1.145 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.32 0.45 0.91 0.54 ;
      RECT 0.82 0.17 0.91 0.54 ;
      RECT 0.32 0.275 0.41 0.54 ;
      RECT 1.38 0.17 1.47 0.4 ;
      RECT 0.82 0.17 1.47 0.26 ;
  END
END OAI32X0P5H7R

MACRO OAI32X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32X0P7H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.335 1.015 1.425 1.48 ;
        RECT 0.07 1.015 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.545 -0.08 0.685 0.385 ;
        RECT 0.07 -0.08 0.16 0.425 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.42 1.055 0.575 1.145 ;
        RECT 0.42 0.71 0.51 1.145 ;
      LAYER MET2 ;
        RECT 0.45 0.84 0.55 1.22 ;
      LAYER VIA1 ;
        RECT 0.455 1.055 0.545 1.145 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.605 0.655 0.805 0.765 ;
        RECT 0.605 0.655 0.695 0.945 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.29 0.625 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.855 0.995 0.945 ;
        RECT 0.905 0.725 0.995 0.945 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.045 0.35 1.215 0.44 ;
        RECT 0.795 1.055 1.175 1.145 ;
        RECT 1.085 0.35 1.175 1.145 ;
      LAYER MET2 ;
        RECT 1.05 0.84 1.15 1.22 ;
      LAYER VIA1 ;
        RECT 1.055 1.055 1.145 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.32 0.475 0.91 0.565 ;
      RECT 0.82 0.17 0.91 0.565 ;
      RECT 0.32 0.3 0.41 0.565 ;
      RECT 1.38 0.17 1.47 0.425 ;
      RECT 0.82 0.17 1.47 0.26 ;
  END
END OAI32X0P7H7R

MACRO OAI32X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32X1H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.355 1.01 1.445 1.48 ;
        RECT 0.07 1.01 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.545 -0.08 0.685 0.35 ;
        RECT 0.07 -0.08 0.16 0.39 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.42 0.62 0.545 0.84 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.675 0.745 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.595 1.405 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.85 0.625 0.985 0.825 ;
      LAYER MET2 ;
        RECT 0.85 0.25 0.95 0.785 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.075 0.35 1.215 0.44 ;
        RECT 0.795 1.05 1.165 1.145 ;
        RECT 1.075 0.35 1.165 1.145 ;
      LAYER MET2 ;
        RECT 0.85 1.015 0.95 1.22 ;
      LAYER VIA1 ;
        RECT 0.855 1.055 0.945 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.32 0.44 0.91 0.53 ;
      RECT 0.82 0.17 0.91 0.53 ;
      RECT 0.32 0.325 0.41 0.53 ;
      RECT 1.355 0.17 1.445 0.39 ;
      RECT 0.82 0.17 1.445 0.26 ;
  END
END OAI32X1H7R

MACRO OAI32X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32X1P4H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.355 1.055 1.445 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 0.545 -0.08 0.685 0.315 ;
        RECT 0.07 -0.08 0.16 0.355 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.62 0.545 0.82 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.675 0.745 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.595 1.405 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.85 0.625 0.985 0.825 ;
      LAYER MET2 ;
        RECT 0.85 0.25 0.95 0.785 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.075 0.35 1.215 0.44 ;
        RECT 0.795 1.055 1.165 1.145 ;
        RECT 1.075 0.35 1.165 1.145 ;
      LAYER MET2 ;
        RECT 0.85 1.015 0.95 1.22 ;
      LAYER VIA1 ;
        RECT 0.855 1.055 0.945 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.32 0.405 0.91 0.495 ;
      RECT 0.82 0.17 0.91 0.495 ;
      RECT 0.32 0.325 0.41 0.495 ;
      RECT 1.355 0.17 1.445 0.355 ;
      RECT 0.82 0.17 1.445 0.26 ;
  END
END OAI32X1P4H7R

MACRO OAI32X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32X2H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.568 1.055 1.658 1.48 ;
        RECT 0.283 1.055 0.373 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 0.783 -0.08 0.873 0.33 ;
        RECT 0.283 -0.08 0.373 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.625 0.435 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.61 0.615 0.745 0.815 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.615 0.958 0.975 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.473 0.655 1.775 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.615 1.203 0.8 ;
      LAYER MET2 ;
        RECT 1.05 0.25 1.15 0.785 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.268 0.35 1.408 0.44 ;
        RECT 1.008 1.055 1.383 1.145 ;
        RECT 1.293 0.35 1.383 1.145 ;
      LAYER MET2 ;
        RECT 1.05 1.015 1.15 1.22 ;
      LAYER VIA1 ;
        RECT 1.055 1.055 1.145 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.533 0.42 1.123 0.51 ;
      RECT 1.033 0.17 1.123 0.51 ;
      RECT 0.533 0.37 0.623 0.51 ;
      RECT 1.568 0.17 1.658 0.345 ;
      RECT 1.033 0.17 1.658 0.26 ;
  END
END OAI32X2H7R

MACRO OAI32X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32X3H7R 0 0 ;
  SIZE 3 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3 1.48 ;
        RECT 2.225 1.24 2.365 1.48 ;
        RECT 0.785 1.24 0.925 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3 0.08 ;
        RECT 1.37 -0.08 1.51 0.175 ;
        RECT 0.84 -0.08 0.98 0.175 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.685 0.455 1.025 0.61 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.7 1.345 0.79 ;
        RECT 1.205 0.66 1.345 0.79 ;
        RECT 0.45 0.625 0.545 0.79 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.17 0.88 1.6 0.97 ;
        RECT 1.51 0.69 1.6 0.97 ;
        RECT 0.17 0.855 0.375 0.97 ;
        RECT 0.17 0.69 0.26 0.97 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.125 0.655 2.465 0.745 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.87 0.835 2.745 0.925 ;
        RECT 2.655 0.625 2.745 0.925 ;
        RECT 1.87 0.69 1.96 0.925 ;
      LAYER MET2 ;
        RECT 2.65 0.43 2.75 0.96 ;
      LAYER VIA1 ;
        RECT 2.655 0.655 2.745 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.045 1.06 2.855 1.15 ;
        RECT 2.475 0.35 2.615 0.44 ;
        RECT 1.69 0.455 2.565 0.565 ;
        RECT 2.475 0.35 2.565 0.565 ;
        RECT 1.945 0.35 2.085 0.565 ;
        RECT 1.69 0.455 1.78 1.15 ;
      LAYER MET2 ;
        RECT 1.85 0.225 1.95 0.76 ;
      LAYER VIA1 ;
        RECT 1.855 0.455 1.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.75 0.17 2.84 0.375 ;
      RECT 0.045 0.275 1.75 0.365 ;
      RECT 1.66 0.17 1.75 0.365 ;
      RECT 2.235 0.17 2.325 0.36 ;
      RECT 1.66 0.17 2.84 0.26 ;
  END
END OAI32X3H7R

MACRO OAI32X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32X4H7R 0 0 ;
  SIZE 5.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.8 1.48 ;
        RECT 4.995 1.225 5.135 1.48 ;
        RECT 4.465 1.225 4.605 1.48 ;
        RECT 0.795 1.03 0.935 1.48 ;
        RECT 0.295 1.03 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.8 0.08 ;
        RECT 3.12 -0.08 3.26 0.26 ;
        RECT 2.59 -0.08 2.73 0.26 ;
        RECT 1.795 -0.08 1.935 0.32 ;
        RECT 1.295 -0.08 1.435 0.32 ;
        RECT 0.795 -0.08 0.935 0.32 ;
        RECT 0.295 -0.08 0.435 0.32 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.245 0.655 0.985 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.245 0.655 1.985 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.56 0.655 3.3 0.745 ;
      LAYER MET2 ;
        RECT 2.85 0.43 2.95 0.96 ;
      LAYER VIA1 ;
        RECT 2.855 0.655 2.945 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.405 0.655 5.145 0.745 ;
      LAYER MET2 ;
        RECT 4.65 0.425 4.75 0.96 ;
      LAYER VIA1 ;
        RECT 4.655 0.655 4.745 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.15 0.835 5.455 0.925 ;
        RECT 5.365 0.74 5.455 0.925 ;
        RECT 4.15 0.655 4.24 0.925 ;
        RECT 3.82 0.655 4.24 0.745 ;
      LAYER MET2 ;
        RECT 3.85 0.43 3.95 0.96 ;
      LAYER VIA1 ;
        RECT 3.855 0.655 3.945 0.745 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.545 1.025 5.745 1.175 ;
        RECT 5.545 0.35 5.635 1.175 ;
        RECT 3.59 0.35 5.635 0.44 ;
        RECT 3.92 0.85 4.06 1.05 ;
        RECT 2.325 0.85 4.06 0.94 ;
        RECT 3.59 0.35 3.68 0.94 ;
        RECT 3.425 0.85 3.515 1.075 ;
        RECT 2.855 0.85 2.995 1.05 ;
        RECT 2.325 0.85 2.465 1.05 ;
      LAYER MET2 ;
        RECT 5.65 0.84 5.75 1.22 ;
      LAYER VIA1 ;
        RECT 5.655 1.055 5.745 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.41 2.16 0.5 ;
      RECT 2.07 0.22 2.16 0.5 ;
      RECT 3.41 0.17 3.5 0.44 ;
      RECT 2.07 0.35 3.5 0.44 ;
      RECT 1.57 0.235 1.66 0.5 ;
      RECT 1.07 0.235 1.16 0.5 ;
      RECT 0.57 0.235 0.66 0.5 ;
      RECT 0.07 0.22 0.16 0.5 ;
      RECT 3.41 0.17 5.665 0.26 ;
      RECT 3.67 1.14 4.29 1.23 ;
      RECT 4.2 1.03 4.29 1.23 ;
      RECT 3.67 1.03 3.81 1.23 ;
      RECT 4.2 1.03 5.4 1.12 ;
      RECT 1.295 1.14 3.245 1.23 ;
      RECT 3.105 1.03 3.245 1.23 ;
      RECT 2.575 1.03 2.715 1.23 ;
      RECT 1.795 1.03 1.935 1.23 ;
      RECT 1.295 1.03 1.435 1.23 ;
      RECT 0.07 0.85 0.16 1.09 ;
      RECT 1.07 0.85 1.16 1.075 ;
      RECT 0.57 0.85 0.66 1.075 ;
      RECT 2.045 0.85 2.185 1.05 ;
      RECT 1.545 0.85 1.685 1.05 ;
      RECT 0.07 0.85 2.185 0.94 ;
  END
END OAI32X4H7R

MACRO OAI33X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33X0P5H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.575 1.225 1.715 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 0.545 -0.08 0.685 0.36 ;
        RECT 0.07 -0.08 0.16 0.4 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.855 0.575 0.945 ;
        RECT 0.425 0.695 0.515 0.945 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.605 0.63 0.805 0.765 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.375 0.63 1.575 0.765 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.195 0.855 1.375 0.945 ;
        RECT 1.195 0.695 1.285 0.945 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.855 1 0.945 ;
        RECT 0.91 0.695 1 0.945 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.81 1.035 1.755 1.125 ;
        RECT 1.665 0.17 1.755 1.125 ;
        RECT 1.56 0.17 1.755 0.375 ;
        RECT 1.06 0.17 1.755 0.26 ;
        RECT 1.06 0.17 1.2 0.36 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.56 ;
      LAYER VIA1 ;
        RECT 1.655 0.255 1.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.32 0.45 1.45 0.54 ;
      RECT 1.31 0.35 1.45 0.54 ;
      RECT 0.835 0.325 0.925 0.54 ;
      RECT 0.32 0.325 0.41 0.54 ;
  END
END OAI33X0P5H7R

MACRO OAI33X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33X0P7H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.575 1.225 1.715 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 0.545 -0.08 0.685 0.36 ;
        RECT 0.07 -0.08 0.16 0.4 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.855 0.575 0.945 ;
        RECT 0.425 0.705 0.515 0.945 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.63 0.825 0.765 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.375 0.63 1.575 0.765 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.185 0.855 1.375 0.945 ;
        RECT 1.185 0.745 1.275 0.945 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.855 1.02 0.945 ;
        RECT 0.93 0.75 1.02 0.945 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.81 1.035 1.755 1.125 ;
        RECT 1.665 0.17 1.755 1.125 ;
        RECT 1.59 0.17 1.755 0.375 ;
        RECT 1.06 0.17 1.755 0.26 ;
        RECT 1.06 0.17 1.2 0.36 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.56 ;
      LAYER VIA1 ;
        RECT 1.655 0.255 1.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.32 0.45 1.465 0.54 ;
      RECT 1.325 0.35 1.465 0.54 ;
      RECT 0.835 0.3 0.925 0.54 ;
      RECT 0.32 0.3 0.41 0.54 ;
  END
END OAI33X0P7H7R

MACRO OAI33X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33X1H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.56 1.225 1.7 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 0.545 -0.08 0.685 0.35 ;
        RECT 0.07 -0.08 0.16 0.39 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.26 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.395 0.625 0.545 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.855 0.79 0.945 ;
        RECT 0.67 0.705 0.76 0.945 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.45 0.625 1.56 0.8 ;
        RECT 1.385 0.625 1.56 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.2 0.855 1.375 0.945 ;
        RECT 1.2 0.73 1.29 0.945 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.85 0.625 1.03 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.795 1.045 1.75 1.135 ;
        RECT 1.65 0.17 1.75 1.135 ;
        RECT 1.6 0.17 1.75 0.365 ;
        RECT 1.045 0.17 1.75 0.26 ;
        RECT 1.045 0.17 1.185 0.35 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.56 ;
      LAYER VIA1 ;
        RECT 1.655 0.255 1.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.32 0.445 1.435 0.535 ;
      RECT 1.295 0.35 1.435 0.535 ;
      RECT 0.82 0.44 1.435 0.535 ;
      RECT 0.32 0.325 0.41 0.535 ;
      RECT 0.82 0.325 0.91 0.535 ;
  END
END OAI33X1H7R

MACRO OAI33X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33X1P4H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.575 1.225 1.715 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 0.545 -0.08 0.685 0.315 ;
        RECT 0.07 -0.08 0.16 0.355 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.855 0.575 0.945 ;
        RECT 0.425 0.661 0.515 0.945 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.605 0.63 0.805 0.765 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.465 0.585 1.565 0.945 ;
        RECT 1.43 0.585 1.565 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.225 0.855 1.375 0.945 ;
        RECT 1.225 0.661 1.315 0.945 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.855 1 0.945 ;
        RECT 0.91 0.661 1 0.945 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.81 1.035 1.745 1.125 ;
        RECT 1.655 0.17 1.745 1.125 ;
        RECT 1.615 0.17 1.745 0.36 ;
        RECT 1.06 0.17 1.745 0.26 ;
        RECT 1.06 0.17 1.2 0.315 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.56 ;
      LAYER VIA1 ;
        RECT 1.655 0.255 1.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.32 0.405 1.465 0.495 ;
      RECT 1.325 0.35 1.465 0.495 ;
      RECT 0.835 0.315 0.925 0.495 ;
      RECT 0.32 0.315 0.41 0.495 ;
  END
END OAI33X1P4H7R

MACRO OAI33X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33X2H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.845 1.055 1.935 1.48 ;
        RECT 0.257 0.88 0.397 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 0.76 -0.08 0.9 0.305 ;
        RECT 0.282 -0.08 0.372 0.345 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.625 0.435 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.615 0.745 0.84 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.615 0.955 0.975 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.63 0.575 1.765 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.425 0.855 1.575 0.945 ;
        RECT 1.425 0.615 1.515 0.945 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.615 1.227 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.665 0.875 1.945 0.965 ;
        RECT 1.855 0.215 1.945 0.965 ;
        RECT 1.805 0.215 1.945 0.32 ;
        RECT 1.274 0.215 1.945 0.305 ;
        RECT 1.022 1.04 1.755 1.13 ;
        RECT 1.665 0.875 1.755 1.13 ;
      LAYER MET2 ;
        RECT 1.85 0.18 1.95 0.56 ;
      LAYER VIA1 ;
        RECT 1.855 0.255 1.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.507 0.395 1.68 0.485 ;
  END
END OAI33X2H7R

MACRO OAI33X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33X3H7R 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.8 1.48 ;
        RECT 3.345 1.095 3.485 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.8 0.08 ;
        RECT 1.54 -0.08 1.68 0.245 ;
        RECT 0.795 -0.08 0.935 0.335 ;
        RECT 0.295 -0.08 0.435 0.335 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.195 0.655 0.535 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.695 0.655 1.035 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.425 0.655 1.765 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.92 0.655 2.265 0.745 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.715 0.655 3.055 0.745 ;
      LAYER MET2 ;
        RECT 2.85 0.43 2.95 0.96 ;
      LAYER VIA1 ;
        RECT 2.855 0.655 2.945 0.745 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.245 0.655 3.585 0.745 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.055 0.425 3.485 0.515 ;
        RECT 3.345 0.35 3.485 0.515 ;
        RECT 2.815 0.35 2.955 0.515 ;
        RECT 2.355 0.735 2.545 0.825 ;
        RECT 2.455 0.425 2.545 0.825 ;
        RECT 2.305 0.915 2.445 1.045 ;
        RECT 2.355 0.735 2.445 1.045 ;
        RECT 1.275 0.915 2.445 1.005 ;
        RECT 2.055 0.35 2.195 0.515 ;
        RECT 1.805 0.915 1.945 1.045 ;
        RECT 1.275 0.915 1.415 1.045 ;
      LAYER MET2 ;
        RECT 2.45 0.425 2.55 0.96 ;
      LAYER VIA1 ;
        RECT 2.455 0.655 2.545 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 3.595 0.915 3.735 1.045 ;
      RECT 3.065 0.915 3.205 1.045 ;
      RECT 2.535 0.915 2.675 1.045 ;
      RECT 2.535 0.915 3.735 1.005 ;
      RECT 0.07 0.425 1.135 0.515 ;
      RECT 1.83 0.17 1.92 0.425 ;
      RECT 1.045 0.335 1.92 0.425 ;
      RECT 0.57 0.31 0.66 0.515 ;
      RECT 0.07 0.295 0.16 0.515 ;
      RECT 3.62 0.17 3.71 0.375 ;
      RECT 3.08 0.17 3.22 0.335 ;
      RECT 2.425 0.17 2.565 0.335 ;
      RECT 1.83 0.17 3.71 0.26 ;
      RECT 2.055 1.14 2.955 1.23 ;
      RECT 2.815 1.095 2.955 1.23 ;
      RECT 2.055 1.095 2.195 1.23 ;
      RECT 0.795 1.14 1.665 1.23 ;
      RECT 1.525 1.095 1.665 1.23 ;
      RECT 0.795 1.095 0.935 1.23 ;
      RECT 0.07 0.915 0.16 1.06 ;
      RECT 1.045 0.915 1.185 1.045 ;
      RECT 0.545 0.915 0.685 1.045 ;
      RECT 0.07 0.915 1.185 1.005 ;
  END
END OAI33X3H7R

MACRO OAI33X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33X4H7R 0 0 ;
  SIZE 4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4 1.48 ;
        RECT 3.425 1.07 3.515 1.48 ;
        RECT 0.465 1.07 0.555 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4 0.08 ;
        RECT 1.64 -0.08 1.78 0.305 ;
        RECT 1.01 -0.08 1.15 0.305 ;
        RECT 0.51 -0.08 0.65 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.37 0.655 0.71 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.87 0.655 1.21 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.54 0.655 1.88 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.04 0.655 2.38 0.745 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.77 0.655 3.11 0.745 ;
      LAYER MET2 ;
        RECT 2.85 0.43 2.95 0.96 ;
      LAYER VIA1 ;
        RECT 2.855 0.655 2.945 0.745 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.26 0.655 3.6 0.745 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.17 0.395 3.47 0.485 ;
        RECT 1.42 0.885 2.56 0.975 ;
        RECT 2.47 0.395 2.56 0.975 ;
        RECT 2.435 0.395 2.56 0.575 ;
      LAYER MET2 ;
        RECT 2.45 0.225 2.55 0.76 ;
      LAYER VIA1 ;
        RECT 2.455 0.455 2.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.285 0.395 2.035 0.485 ;
      RECT 1.945 0.215 2.035 0.485 ;
      RECT 0.285 0.33 0.375 0.485 ;
      RECT 3.605 0.215 3.695 0.355 ;
      RECT 1.945 0.215 3.695 0.305 ;
      RECT 2.65 0.885 3.79 0.975 ;
      RECT 2.17 1.095 3.04 1.185 ;
      RECT 0.94 1.095 1.81 1.185 ;
      RECT 0.19 0.885 1.33 0.975 ;
  END
END OAI33X4H7R

MACRO OAO211X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAO211X0P5H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.505 1.04 1.595 1.48 ;
        RECT 0.77 1.205 0.91 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.36 -0.08 1.45 0.37 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.615 0.545 0.84 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.455 0.895 0.555 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.005 0.625 1.185 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.755 0.255 1.845 1.14 ;
        RECT 1.595 0.255 1.845 0.36 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.56 ;
      LAYER VIA1 ;
        RECT 1.655 0.255 1.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.275 0.485 1.365 1.14 ;
      RECT 1.275 0.64 1.665 0.73 ;
      RECT 1.235 0.397 1.275 0.525 ;
      RECT 1.235 0.44 1.321 0.525 ;
      RECT 1.189 0.354 1.235 0.482 ;
      RECT 1.143 0.308 1.189 0.436 ;
      RECT 1.105 0.354 1.235 0.394 ;
      RECT 1 0.285 1.143 0.375 ;
      RECT 0.505 1.025 1.14 1.115 ;
      RECT 0.045 0.27 0.715 0.36 ;
  END
END OAO211X0P5H7R

MACRO OAO211X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAO211X0P7H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.49 1.04 1.58 1.48 ;
        RECT 0.755 1.06 0.895 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.345 -0.08 1.435 0.37 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.365 0.625 0.545 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.45 0.85 0.57 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.99 0.625 1.17 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.74 0.255 1.83 1.108 ;
        RECT 1.58 0.255 1.83 0.36 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.56 ;
      LAYER VIA1 ;
        RECT 1.655 0.255 1.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.26 0.485 1.35 1.14 ;
      RECT 1.26 0.64 1.65 0.73 ;
      RECT 1.22 0.397 1.26 0.525 ;
      RECT 1.22 0.44 1.306 0.525 ;
      RECT 1.174 0.354 1.22 0.482 ;
      RECT 1.128 0.308 1.174 0.436 ;
      RECT 1.09 0.354 1.22 0.394 ;
      RECT 0.985 0.285 1.128 0.375 ;
      RECT 1.01 0.88 1.1 1.145 ;
      RECT 0.53 0.88 0.62 1.12 ;
      RECT 0.53 0.88 1.1 0.97 ;
      RECT 0.045 0.27 0.715 0.36 ;
  END
END OAO211X0P7H7R

MACRO OAO211X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAO211X1H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.49 1.055 1.58 1.48 ;
        RECT 0.755 1.06 0.895 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.35 -0.08 1.44 0.37 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.365 0.625 0.545 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.45 0.85 0.57 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.99 0.625 1.17 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.74 0.255 1.83 1.075 ;
        RECT 1.58 0.255 1.83 0.36 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.56 ;
      LAYER VIA1 ;
        RECT 1.655 0.255 1.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.26 0.48 1.35 1.14 ;
      RECT 1.26 0.64 1.65 0.73 ;
      RECT 1.225 0.394 1.26 0.523 ;
      RECT 1.179 0.354 1.225 0.482 ;
      RECT 1.179 0.435 1.306 0.482 ;
      RECT 1.133 0.308 1.179 0.436 ;
      RECT 1.095 0.285 1.133 0.394 ;
      RECT 0.985 0.285 1.133 0.375 ;
      RECT 1.01 0.88 1.1 1.14 ;
      RECT 0.53 0.88 0.62 1.12 ;
      RECT 0.53 0.88 1.1 0.97 ;
      RECT 0.045 0.27 0.715 0.36 ;
  END
END OAO211X1H7R

MACRO OAO211X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAO211X1P4H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.49 1.055 1.58 1.48 ;
        RECT 0.755 1.06 0.895 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.35 -0.08 1.44 0.37 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.365 0.625 0.545 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.45 0.85 0.57 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.99 0.625 1.17 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.74 0.255 1.83 1.031 ;
        RECT 1.58 0.255 1.83 0.345 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.56 ;
      LAYER VIA1 ;
        RECT 1.655 0.255 1.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.26 0.48 1.35 1.14 ;
      RECT 1.26 0.64 1.65 0.73 ;
      RECT 1.225 0.394 1.26 0.523 ;
      RECT 1.179 0.354 1.225 0.482 ;
      RECT 1.179 0.435 1.306 0.482 ;
      RECT 1.133 0.308 1.179 0.436 ;
      RECT 1.095 0.285 1.133 0.394 ;
      RECT 0.985 0.285 1.133 0.375 ;
      RECT 1.01 0.88 1.1 1.14 ;
      RECT 0.53 0.88 0.62 1.12 ;
      RECT 0.53 0.88 1.1 0.97 ;
      RECT 0.045 0.27 0.715 0.36 ;
  END
END OAO211X1P4H7R

MACRO OAO211X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAO211X2H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.49 1.055 1.58 1.48 ;
        RECT 0.755 1.06 0.895 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.305 -0.08 1.395 0.37 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.365 0.625 0.545 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.62 0.45 0.845 0.57 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.99 0.625 1.17 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.74 0.255 1.83 0.965 ;
        RECT 1.53 0.255 1.83 0.345 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.56 ;
      LAYER VIA1 ;
        RECT 1.655 0.255 1.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.26 0.525 1.35 1.14 ;
      RECT 1.26 0.64 1.6 0.73 ;
      RECT 1.226 0.44 1.26 0.568 ;
      RECT 1.18 0.4 1.226 0.528 ;
      RECT 1.18 0.48 1.306 0.528 ;
      RECT 1.134 0.354 1.18 0.482 ;
      RECT 1.088 0.308 1.134 0.436 ;
      RECT 1.05 0.354 1.18 0.394 ;
      RECT 0.945 0.285 1.088 0.375 ;
      RECT 1.01 0.88 1.1 1.14 ;
      RECT 0.53 0.88 0.62 1.12 ;
      RECT 0.53 0.88 1.1 0.97 ;
      RECT 0.045 0.27 0.715 0.36 ;
  END
END OAO211X2H7R

MACRO OAO211X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAO211X3H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 2.03 1.055 2.12 1.48 ;
        RECT 1.53 1.055 1.62 1.48 ;
        RECT 0.795 1.06 0.935 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.96 -0.08 2.05 0.37 ;
        RECT 1.345 -0.08 1.435 0.37 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.365 0.625 0.545 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.7 0.455 0.79 0.675 ;
        RECT 0.62 0.455 0.79 0.545 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.03 0.625 1.21 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.78 0.255 1.87 1.045 ;
        RECT 1.625 0.255 1.87 0.345 ;
      LAYER MET2 ;
        RECT 1.65 0.18 1.75 0.56 ;
      LAYER VIA1 ;
        RECT 1.655 0.255 1.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.3 0.525 1.39 1.06 ;
      RECT 1.3 0.64 1.69 0.73 ;
      RECT 1.28 0.447 1.3 0.575 ;
      RECT 1.234 0.414 1.28 0.542 ;
      RECT 1.234 0.48 1.346 0.542 ;
      RECT 1.188 0.368 1.234 0.496 ;
      RECT 1.15 0.345 1.188 0.454 ;
      RECT 1.025 0.345 1.188 0.435 ;
      RECT 1.05 0.88 1.14 1.06 ;
      RECT 0.57 0.88 0.66 1.04 ;
      RECT 0.57 0.88 1.14 0.97 ;
      RECT 0.045 0.27 0.715 0.36 ;
  END
END OAO211X3H7R

MACRO OAO211X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAO211X4H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 2.09 1.055 2.18 1.48 ;
        RECT 1.59 1.055 1.68 1.48 ;
        RECT 0.855 1.08 0.995 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 2.005 -0.08 2.095 0.345 ;
        RECT 1.34 -0.08 1.43 0.33 ;
        RECT 0.36 -0.08 0.5 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.43 0.625 0.61 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.8 0.455 0.975 0.545 ;
        RECT 0.8 0.455 0.89 0.67 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1 0.655 1.27 0.755 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.84 0.825 1.97 0.975 ;
        RECT 1.84 0.395 1.93 0.975 ;
        RECT 1.68 0.395 1.93 0.485 ;
      LAYER MET2 ;
        RECT 1.85 0.625 1.95 1.16 ;
      LAYER VIA1 ;
        RECT 1.855 0.855 1.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.36 0.55 1.45 1.035 ;
      RECT 1.36 0.64 1.75 0.73 ;
      RECT 1.347 0.475 1.36 0.604 ;
      RECT 1.301 0.446 1.347 0.574 ;
      RECT 1.301 0.505 1.406 0.574 ;
      RECT 1.255 0.4 1.301 0.528 ;
      RECT 1.209 0.354 1.255 0.482 ;
      RECT 1.163 0.308 1.209 0.436 ;
      RECT 1.125 0.354 1.255 0.394 ;
      RECT 1.02 0.285 1.163 0.375 ;
      RECT 1.11 0.9 1.2 1.04 ;
      RECT 0.605 0.9 0.745 0.995 ;
      RECT 0.605 0.9 1.2 0.99 ;
      RECT 0.045 0.27 0.815 0.36 ;
  END
END OAO211X4H7R

MACRO OAOI211X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAOI211X0P5H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.79 1.205 0.93 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.346 -0.08 1.436 0.37 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 0.625 0.55 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.7 0.455 0.79 0.68 ;
        RECT 0.625 0.455 0.79 0.545 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.635 1.22 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.6 1.15 1.135 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.315 0.535 1.405 1.14 ;
        RECT 1.267 0.49 1.361 0.57 ;
        RECT 1.221 0.466 1.315 0.524 ;
        RECT 1.313 0.535 1.405 0.594 ;
        RECT 1.175 0.442 1.313 0.478 ;
        RECT 1.157 0.396 1.267 0.446 ;
        RECT 1.111 0.35 1.221 0.414 ;
        RECT 1.065 0.255 1.175 0.368 ;
        RECT 1.022 0.255 1.175 0.345 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.385 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.525 1.025 1.18 1.115 ;
      RECT 0.045 0.27 0.715 0.36 ;
  END
END OAOI211X0P5H7R

MACRO OAOI211X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAOI211X0P7H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.79 1.173 0.93 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.306 -0.08 1.396 0.37 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 0.625 0.55 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.7 0.455 0.79 0.675 ;
        RECT 0.62 0.455 0.79 0.545 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.98 0.655 1.205 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.6 1.15 1.135 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.295 0.555 1.385 1.108 ;
        RECT 1.221 0.51 1.341 0.564 ;
        RECT 1.175 0.473 1.295 0.518 ;
        RECT 1.267 0.555 1.385 0.601 ;
        RECT 1.163 0.436 1.267 0.489 ;
        RECT 1.117 0.39 1.221 0.46 ;
        RECT 1.071 0.255 1.175 0.414 ;
        RECT 1.025 0.255 1.175 0.368 ;
        RECT 1.02 0.255 1.175 0.345 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.385 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.525 0.993 1.16 1.083 ;
      RECT 0.045 0.27 0.715 0.36 ;
  END
END OAOI211X0P7H7R

MACRO OAOI211X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAOI211X1H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.79 1.125 0.93 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.336 -0.08 1.426 0.37 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.625 0.545 0.825 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.7 0.455 0.79 0.68 ;
        RECT 0.625 0.455 0.79 0.545 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.625 1.205 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.6 1.15 1.135 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.295 0.525 1.385 1.06 ;
        RECT 1.221 0.48 1.341 0.534 ;
        RECT 1.175 0.443 1.295 0.488 ;
        RECT 1.267 0.525 1.385 0.571 ;
        RECT 1.147 0.406 1.267 0.451 ;
        RECT 1.101 0.36 1.221 0.414 ;
        RECT 1.055 0.255 1.175 0.368 ;
        RECT 1.02 0.255 1.175 0.345 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.385 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.525 0.945 1.16 1.035 ;
      RECT 0.045 0.27 0.715 0.36 ;
  END
END OAOI211X1H7R

MACRO OAOI211X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAOI211X1P4H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 0.875 1.08 1.015 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.385 -0.08 1.475 0.345 ;
        RECT 0.36 -0.08 0.5 0.175 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.395 0.645 0.665 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.26 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.8 0.455 0.975 0.545 ;
        RECT 0.8 0.455 0.89 0.67 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.02 0.655 1.29 0.755 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.38 0.825 1.545 1.031 ;
        RECT 1.38 0.54 1.47 1.031 ;
        RECT 1.34 0.495 1.426 0.58 ;
        RECT 1.294 0.452 1.38 0.537 ;
        RECT 1.248 0.409 1.34 0.491 ;
        RECT 1.102 0.363 1.294 0.43 ;
        RECT 1.102 0.34 1.248 0.43 ;
        RECT 1.21 0.409 1.34 0.449 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.13 0.9 1.22 1.04 ;
      RECT 0.625 0.9 0.765 1.03 ;
      RECT 0.625 0.9 1.22 0.99 ;
      RECT 0.045 0.27 0.815 0.36 ;
  END
END OAOI211X1P4H7R

MACRO OAOI211X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAOI211X2H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 0.995 1.055 1.085 1.48 ;
        RECT 0.285 1.055 0.375 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.425 -0.08 1.515 0.345 ;
        RECT 0.51 -0.08 0.65 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.595 0.615 0.775 0.765 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.625 0.435 0.775 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.88 0.655 1.18 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.355 0.625 1.548 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.45 0.885 1.745 0.975 ;
        RECT 1.655 0.445 1.745 0.975 ;
        RECT 1.175 0.445 1.745 0.535 ;
        RECT 1.175 0.37 1.265 0.535 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.285 0.395 0.9 0.485 ;
      RECT 0.285 0.32 0.375 0.485 ;
      RECT 0.72 0.875 1.34 0.965 ;
  END
END OAOI211X2H7R

MACRO OAOI211X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAOI211X3H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 1.525 1.095 1.665 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 2.055 -0.08 2.195 0.305 ;
        RECT 0.795 -0.08 0.935 0.335 ;
        RECT 0.295 -0.08 0.435 0.335 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.665 0.655 1.005 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.165 0.655 0.505 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.195 0.655 1.735 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.9 0.655 2.24 0.745 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.025 0.855 2.42 0.945 ;
        RECT 2.33 0.28 2.42 0.945 ;
        RECT 1.31 0.44 2.42 0.53 ;
        RECT 1.805 0.41 2.42 0.53 ;
        RECT 2.025 0.855 2.165 1.02 ;
        RECT 1.805 0.305 1.945 0.53 ;
        RECT 1.31 0.35 1.45 0.53 ;
      LAYER MET2 ;
        RECT 2.25 0.63 2.35 1.16 ;
      LAYER VIA1 ;
        RECT 2.255 0.855 2.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.8 1.11 2.39 1.2 ;
      RECT 2.3 1.055 2.39 1.2 ;
      RECT 1.8 0.9 1.89 1.2 ;
      RECT 1.275 0.9 1.415 1.035 ;
      RECT 0.795 0.9 0.935 1.02 ;
      RECT 0.795 0.9 1.89 0.99 ;
      RECT 0.07 0.425 1.16 0.515 ;
      RECT 1.07 0.17 1.16 0.515 ;
      RECT 0.57 0.28 0.66 0.515 ;
      RECT 0.07 0.28 0.16 0.515 ;
      RECT 1.575 0.17 1.715 0.35 ;
      RECT 1.07 0.17 1.715 0.26 ;
      RECT 0.57 1.11 1.185 1.2 ;
      RECT 1.045 1.08 1.185 1.2 ;
      RECT 0.57 0.915 0.66 1.2 ;
      RECT 0.07 0.915 0.16 1.06 ;
      RECT 0.07 0.915 0.66 1.005 ;
  END
END OAOI211X3H7R

MACRO OAOI211X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAOI211X4H7R 0 0 ;
  SIZE 3 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3 1.48 ;
        RECT 1.737 1.095 1.877 1.48 ;
        RECT 0.507 1.095 0.647 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3 0.08 ;
        RECT 2.267 -0.08 2.407 0.305 ;
        RECT 1.007 -0.08 1.147 0.305 ;
        RECT 0.507 -0.08 0.647 0.305 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.877 0.655 1.217 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.377 0.655 0.717 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.407 0.655 1.947 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.112 0.655 2.452 0.745 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.237 0.855 2.632 0.945 ;
        RECT 2.542 0.325 2.632 0.945 ;
        RECT 1.522 0.41 2.632 0.5 ;
        RECT 2.237 0.855 2.377 0.975 ;
        RECT 2.017 0.38 2.157 0.5 ;
        RECT 1.522 0.395 1.662 0.5 ;
      LAYER MET2 ;
        RECT 2.45 0.625 2.55 1.16 ;
      LAYER VIA1 ;
        RECT 2.455 0.855 2.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.012 1.065 2.627 1.155 ;
      RECT 2.012 0.9 2.102 1.155 ;
      RECT 1.007 0.9 2.102 0.99 ;
      RECT 0.282 0.395 1.372 0.485 ;
      RECT 1.282 0.17 1.372 0.485 ;
      RECT 0.282 0.31 0.372 0.485 ;
      RECT 1.787 0.17 1.927 0.32 ;
      RECT 1.282 0.17 1.927 0.26 ;
      RECT 0.782 1.08 1.397 1.17 ;
      RECT 0.782 0.915 0.872 1.17 ;
      RECT 0.257 0.915 0.872 1.005 ;
  END
END OAOI211X4H7R

MACRO OR2X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X0P5H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.555 1.005 0.695 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.555 -0.08 0.695 0.325 ;
        RECT 0.045 -0.08 0.185 0.34 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.625 0.57 0.86 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.69 0.345 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.84 0.225 0.945 1.085 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.56 ;
      LAYER VIA1 ;
        RECT 0.855 0.255 0.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.43 0.16 1.075 ;
      RECT 0.66 0.43 0.75 0.575 ;
      RECT 0.07 0.43 0.75 0.52 ;
      RECT 0.32 0.215 0.41 0.52 ;
  END
END OR2X0P5H7R

MACRO OR2X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X0P7H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.58 0.975 0.67 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.58 -0.08 0.67 0.33 ;
        RECT 0.045 -0.08 0.185 0.32 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.625 0.57 0.85 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.69 0.345 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.805 0.945 0.945 1.035 ;
        RECT 0.855 0.23 0.945 1.035 ;
        RECT 0.805 0.23 0.945 0.32 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.445 0.16 1.06 ;
      RECT 0.675 0.445 0.765 0.585 ;
      RECT 0.07 0.445 0.765 0.535 ;
      RECT 0.32 0.22 0.41 0.535 ;
  END
END OR2X0P7H7R

MACRO OR2X12H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X12H7R 0 0 ;
  SIZE 3.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.4 1.48 ;
        RECT 3.067 1.055 3.157 1.48 ;
        RECT 2.567 1.07 2.657 1.48 ;
        RECT 2.067 1.07 2.157 1.48 ;
        RECT 1.567 1.055 1.657 1.48 ;
        RECT 0.572 1.07 0.662 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.4 0.08 ;
        RECT 3.028 -0.08 3.118 0.345 ;
        RECT 2.503 -0.08 2.643 0.305 ;
        RECT 2.003 -0.08 2.143 0.305 ;
        RECT 1.297 -0.08 1.437 0.305 ;
        RECT 0.797 -0.08 0.937 0.305 ;
        RECT 0.322 -0.08 0.412 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.417 0.655 0.757 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.917 0.655 1.257 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.792 0.855 2.932 0.945 ;
        RECT 2.842 0.395 2.932 0.945 ;
        RECT 1.753 0.395 2.932 0.485 ;
      LAYER MET2 ;
        RECT 2.65 0.63 2.75 1.16 ;
      LAYER VIA1 ;
        RECT 2.655 0.855 2.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.047 0.885 1.437 0.975 ;
      RECT 1.347 0.395 1.437 0.975 ;
      RECT 1.347 0.625 2.752 0.715 ;
      RECT 0.547 0.395 1.437 0.485 ;
      RECT 0.847 1.065 1.437 1.155 ;
      RECT 0.847 0.865 0.937 1.155 ;
      RECT 0.297 0.865 0.937 0.955 ;
  END
END OR2X12H7R

MACRO OR2X16H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X16H7R 0 0 ;
  SIZE 4.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.4 1.48 ;
        RECT 4.052 1.055 4.142 1.48 ;
        RECT 3.552 1.07 3.642 1.48 ;
        RECT 3.052 1.07 3.142 1.48 ;
        RECT 2.552 1.07 2.642 1.48 ;
        RECT 2.052 1.055 2.142 1.48 ;
        RECT 0.822 1.07 0.912 1.48 ;
        RECT 0.322 1.055 0.412 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.4 0.08 ;
        RECT 4.028 -0.08 4.118 0.345 ;
        RECT 3.503 -0.08 3.643 0.305 ;
        RECT 3.003 -0.08 3.143 0.305 ;
        RECT 2.503 -0.08 2.643 0.305 ;
        RECT 1.797 -0.08 1.937 0.305 ;
        RECT 1.297 -0.08 1.437 0.305 ;
        RECT 0.797 -0.08 0.937 0.305 ;
        RECT 0.322 -0.08 0.412 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.477 0.655 1.017 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.217 0.655 1.757 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.277 0.855 3.917 0.945 ;
        RECT 3.827 0.395 3.917 0.945 ;
        RECT 2.253 0.395 3.917 0.485 ;
      LAYER MET2 ;
        RECT 3.65 0.63 3.75 1.16 ;
      LAYER VIA1 ;
        RECT 3.655 0.855 3.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.297 0.885 1.937 0.975 ;
      RECT 1.847 0.395 1.937 0.975 ;
      RECT 1.847 0.625 3.707 0.715 ;
      RECT 0.547 0.395 1.937 0.485 ;
      RECT 1.097 1.065 1.687 1.155 ;
      RECT 1.097 0.89 1.187 1.155 ;
      RECT 0.547 0.89 1.187 0.98 ;
  END
END OR2X16H7R

MACRO OR2X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X1H7R 0 0 ;
  SIZE 1.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.2 1.48 ;
        RECT 0.58 0.955 0.67 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.2 0.08 ;
        RECT 0.555 -0.08 0.695 0.34 ;
        RECT 0.045 -0.08 0.185 0.34 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.61 0.57 0.845 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.69 0.345 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.885 0.24 0.975 1.1 ;
        RECT 0.825 0.24 0.975 0.345 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.56 ;
      LAYER VIA1 ;
        RECT 0.855 0.255 0.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.43 0.16 1.095 ;
      RECT 0.705 0.43 0.795 0.635 ;
      RECT 0.07 0.43 0.795 0.52 ;
      RECT 0.295 0.25 0.435 0.52 ;
  END
END OR2X1H7R

MACRO OR2X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X1P4H7R 0 0 ;
  SIZE 1 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1 1.48 ;
        RECT 0.57 1.07 0.66 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1 0.08 ;
        RECT 0.57 -0.08 0.66 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.625 0.56 0.85 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.75 0.345 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.81 0.825 0.955 1.006 ;
        RECT 0.865 0.265 0.955 1.006 ;
        RECT 0.81 0.265 0.955 0.355 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 1.065 0.185 1.155 ;
      RECT 0.045 0.445 0.135 1.155 ;
      RECT 0.685 0.445 0.775 0.651 ;
      RECT 0.045 0.445 0.775 0.535 ;
      RECT 0.32 0.22 0.41 0.535 ;
  END
END OR2X1P4H7R

MACRO OR2X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X2H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.215 0.955 1.305 1.48 ;
        RECT 0.57 1.225 0.71 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.215 -0.08 1.305 0.45 ;
        RECT 0.57 -0.08 0.71 0.425 ;
        RECT 0.07 -0.08 0.16 0.45 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.745 0.6 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.72 0.345 1.175 ;
      LAYER MET2 ;
        RECT 0.25 0.84 0.35 1.22 ;
      LAYER VIA1 ;
        RECT 0.255 1.055 0.345 1.145 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 1.055 1.035 1.145 ;
        RECT 0.945 0.31 1.035 1.145 ;
      LAYER MET2 ;
        RECT 0.85 0.84 0.95 1.22 ;
      LAYER VIA1 ;
        RECT 0.855 1.055 0.945 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.54 0.16 1.08 ;
      RECT 0.07 0.54 0.855 0.63 ;
      RECT 0.32 0.31 0.41 0.63 ;
  END
END OR2X2H7R

MACRO OR2X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X3H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 1.12 1.055 1.21 1.48 ;
        RECT 0.58 1.07 0.67 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 1.12 -0.08 1.21 0.345 ;
        RECT 0.58 -0.08 0.67 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.625 0.575 0.85 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.72 0.35 0.99 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.87 0.225 0.96 1.045 ;
        RECT 0.84 0.225 0.96 0.375 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.56 ;
      LAYER VIA1 ;
        RECT 0.855 0.255 0.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.445 0.16 1.08 ;
      RECT 0.69 0.445 0.78 0.605 ;
      RECT 0.07 0.445 0.78 0.535 ;
      RECT 0.32 0.28 0.41 0.535 ;
  END
END OR2X3H7R

MACRO OR2X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X4H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.305 1.205 1.445 1.48 ;
        RECT 0.775 1.205 0.915 1.48 ;
        RECT 0.07 0.94 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.305 -0.08 1.445 0.175 ;
        RECT 0.79 -0.08 0.93 0.34 ;
        RECT 0.57 -0.08 0.66 0.33 ;
        RECT 0.07 -0.08 0.16 0.353 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.62 0.255 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.62 0.615 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.04 0.805 1.745 0.896 ;
        RECT 1.655 0.265 1.745 0.896 ;
        RECT 1.04 0.265 1.745 0.355 ;
      LAYER MET2 ;
        RECT 1.65 0.23 1.75 0.76 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.545 0.915 0.795 1.005 ;
      RECT 0.705 0.43 0.795 1.005 ;
      RECT 0.705 0.54 1.44 0.63 ;
      RECT 0.32 0.43 0.795 0.52 ;
      RECT 0.32 0.32 0.41 0.52 ;
  END
END OR2X4H7R

MACRO OR2X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X6H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.552 1.07 1.642 1.48 ;
        RECT 1.052 1.055 1.142 1.48 ;
        RECT 0.322 1.055 0.412 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.527 -0.08 1.667 0.305 ;
        RECT 1.052 -0.08 1.142 0.345 ;
        RECT 0.822 -0.08 0.912 0.345 ;
        RECT 0.322 -0.08 0.412 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.645 0.495 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.59 0.615 0.79 0.75 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.277 0.855 1.917 0.945 ;
        RECT 1.827 0.395 1.917 0.945 ;
        RECT 1.802 0.205 1.892 0.485 ;
        RECT 1.277 0.395 1.917 0.485 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.797 0.85 0.97 0.94 ;
      RECT 0.88 0.435 0.97 0.94 ;
      RECT 0.88 0.625 1.692 0.715 ;
      RECT 0.572 0.435 0.97 0.525 ;
      RECT 0.572 0.37 0.662 0.525 ;
  END
END OR2X6H7R

MACRO OR2X8H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X8H7R 0 0 ;
  SIZE 2.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.8 1.48 ;
        RECT 2.33 1.055 2.42 1.48 ;
        RECT 1.83 1.07 1.92 1.48 ;
        RECT 1.33 1.055 1.42 1.48 ;
        RECT 0.31 1.095 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.8 0.08 ;
        RECT 2.33 -0.08 2.42 0.345 ;
        RECT 1.805 -0.08 1.945 0.305 ;
        RECT 1.33 -0.08 1.42 0.345 ;
        RECT 1.06 -0.08 1.2 0.32 ;
        RECT 0.56 -0.08 0.7 0.305 ;
        RECT 0.085 -0.08 0.175 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.18 0.655 0.52 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.68 0.655 1.02 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.555 0.855 2.195 0.945 ;
        RECT 2.105 0.395 2.195 0.945 ;
        RECT 1.555 0.395 2.195 0.485 ;
      LAYER MET2 ;
        RECT 2.05 0.63 2.15 1.16 ;
      LAYER VIA1 ;
        RECT 2.055 0.855 2.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.81 0.905 1.2 0.995 ;
      RECT 1.11 0.41 1.2 0.995 ;
      RECT 1.11 0.625 2.015 0.715 ;
      RECT 0.335 0.41 1.2 0.5 ;
      RECT 0.835 0.32 0.925 0.5 ;
      RECT 0.335 0.32 0.425 0.5 ;
      RECT 0.61 1.085 1.2 1.175 ;
      RECT 0.61 0.905 0.7 1.175 ;
      RECT 0.06 0.905 0.7 0.995 ;
  END
END OR2X8H7R

MACRO OR3X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X0P5H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.915 0.995 1.005 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.9 -0.08 0.99 0.35 ;
        RECT 0.4 -0.08 0.49 0.35 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.82 0.625 0.945 0.845 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.625 0.59 0.825 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.73 0.35 1 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.21 0.225 1.345 1.08 ;
      LAYER MET2 ;
        RECT 1.25 0.18 1.35 0.56 ;
      LAYER VIA1 ;
        RECT 1.255 0.255 1.345 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.44 0.16 1.08 ;
      RECT 1.03 0.44 1.12 0.58 ;
      RECT 0.07 0.44 1.12 0.53 ;
      RECT 0.65 0.24 0.74 0.53 ;
      RECT 0.15 0.225 0.24 0.53 ;
  END
END OR3X0P5H7R

MACRO OR3X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X0P7H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.915 0.995 1.005 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.9 -0.08 0.99 0.35 ;
        RECT 0.4 -0.08 0.49 0.35 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.625 0.835 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.725 0.565 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.245 0.62 0.345 0.89 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.18 0.225 1.345 1.048 ;
      LAYER MET2 ;
        RECT 1.22 0.18 1.32 0.56 ;
      LAYER VIA1 ;
        RECT 1.225 0.255 1.315 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.065 0.98 0.26 1.07 ;
      RECT 0.065 0.44 0.155 1.07 ;
      RECT 1 0.44 1.09 0.599 ;
      RECT 0.065 0.44 1.09 0.53 ;
      RECT 0.65 0.24 0.74 0.53 ;
      RECT 0.145 0.225 0.235 0.53 ;
  END
END OR3X0P7H7R

MACRO OR3X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X1H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.89 1.08 1.03 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.875 -0.08 1.015 0.325 ;
        RECT 0.375 -0.08 0.515 0.325 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.8 0.73 0.945 0.975 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.595 0.595 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.69 0.345 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.21 0.235 1.345 1.13 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.225 0.16 1.17 ;
      RECT 1.03 0.415 1.12 0.665 ;
      RECT 0.07 0.415 1.12 0.505 ;
      RECT 0.625 0.25 0.765 0.505 ;
  END
END OR3X1H7R

MACRO OR3X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X1P4H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.915 0.995 1.005 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.9 -0.08 0.99 0.339 ;
        RECT 0.4 -0.08 0.49 0.339 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.795 0.625 0.945 0.805 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.625 0.595 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.705 0.35 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.215 0.31 1.345 0.975 ;
      LAYER MET2 ;
        RECT 1.25 0.63 1.35 1.16 ;
      LAYER VIA1 ;
        RECT 1.255 0.855 1.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.214 0.16 1.08 ;
      RECT 1.035 0.445 1.125 0.665 ;
      RECT 0.07 0.445 1.125 0.535 ;
      RECT 0.65 0.229 0.74 0.535 ;
  END
END OR3X1P4H7R

MACRO OR3X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X2H7R 0 0 ;
  SIZE 1.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.8 1.48 ;
        RECT 1.46 1.04 1.55 1.48 ;
        RECT 0.94 1.07 1.03 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.8 0.08 ;
        RECT 1.46 -0.08 1.55 0.45 ;
        RECT 0.945 -0.08 1.035 0.24 ;
        RECT 0.415 -0.08 0.505 0.245 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.755 0.83 0.99 0.945 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.75 0.575 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.565 0.35 0.835 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.21 0.3 1.345 1.18 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.335 0.16 1.165 ;
      RECT 1.01 0.335 1.1 0.675 ;
      RECT 0.07 0.335 1.1 0.425 ;
  END
END OR3X2H7R

MACRO OR3X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X3H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.435 0.98 1.525 1.48 ;
        RECT 0.915 0.995 1.005 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.435 -0.08 1.525 0.354 ;
        RECT 0.9 -0.08 0.99 0.339 ;
        RECT 0.4 -0.08 0.49 0.339 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.795 0.625 0.945 0.805 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.625 0.595 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.65 0.345 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.155 0.855 1.345 0.945 ;
        RECT 1.255 0.265 1.345 0.945 ;
        RECT 1.155 0.265 1.345 0.355 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.075 0.274 0.165 1 ;
      RECT 1.075 0.445 1.165 0.665 ;
      RECT 0.075 0.445 1.165 0.535 ;
      RECT 0.65 0.289 0.74 0.535 ;
  END
END OR3X3H7R

MACRO OR3X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X4H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.641 1.06 1.781 1.48 ;
        RECT 0.89 1.06 1.03 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.641 -0.08 1.781 0.34 ;
        RECT 1.12 -0.08 1.26 0.325 ;
        RECT 0.875 -0.08 1.015 0.325 ;
        RECT 0.375 -0.08 0.515 0.325 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.795 0.625 0.945 0.805 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.445 0.595 0.595 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.665 0.345 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.921 0.88 2.145 1.15 ;
        RECT 2.055 0.46 2.145 1.15 ;
        RECT 1.921 0.245 2.061 0.55 ;
        RECT 1.376 0.88 2.145 0.97 ;
        RECT 1.376 0.46 2.145 0.55 ;
        RECT 1.376 0.88 1.516 1.135 ;
        RECT 1.376 0.265 1.516 0.55 ;
      LAYER MET2 ;
        RECT 2.05 0.63 2.15 1.16 ;
      LAYER VIA1 ;
        RECT 2.055 0.855 2.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.31 0.16 1.08 ;
      RECT 1.069 0.665 1.796 0.755 ;
      RECT 1.069 0.415 1.159 0.755 ;
      RECT 0.07 0.415 1.159 0.505 ;
      RECT 0.65 0.31 0.74 0.505 ;
  END
END OR3X4H7R

MACRO OR3X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X6H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.572 1.07 1.662 1.48 ;
        RECT 1.072 1.07 1.162 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.547 -0.08 1.687 0.305 ;
        RECT 1.047 -0.08 1.187 0.305 ;
        RECT 0.547 -0.08 0.687 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.855 0.595 1.005 0.775 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.615 0.745 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.422 0.575 0.557 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.297 0.855 1.937 0.945 ;
        RECT 1.847 0.395 1.937 0.945 ;
        RECT 1.822 0.315 1.912 0.485 ;
        RECT 1.297 0.395 1.937 0.485 ;
      LAYER MET2 ;
        RECT 1.65 0.63 1.75 1.16 ;
      LAYER VIA1 ;
        RECT 1.655 0.855 1.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.242 0.865 0.437 0.955 ;
      RECT 0.242 0.355 0.332 0.955 ;
      RECT 1.107 0.625 1.757 0.715 ;
      RECT 1.107 0.395 1.197 0.715 ;
      RECT 0.242 0.395 1.197 0.485 ;
      RECT 0.242 0.355 0.437 0.485 ;
  END
END OR3X6H7R

MACRO OR3X8H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X8H7R 0 0 ;
  SIZE 3.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.2 1.48 ;
        RECT 2.815 1.055 2.905 1.48 ;
        RECT 2.315 1.07 2.405 1.48 ;
        RECT 1.815 1.07 1.905 1.48 ;
        RECT 1.29 1.08 1.43 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.2 0.08 ;
        RECT 2.815 -0.08 2.905 0.345 ;
        RECT 2.29 -0.08 2.43 0.305 ;
        RECT 1.79 -0.08 1.93 0.305 ;
        RECT 1.29 -0.08 1.43 0.305 ;
        RECT 0.56 -0.08 0.7 0.305 ;
        RECT 0.06 -0.08 0.2 0.32 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.4 0.655 1.74 0.745 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.705 0.655 1.045 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.63 0.53 0.77 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.04 0.855 2.68 0.945 ;
        RECT 2.59 0.395 2.68 0.945 ;
        RECT 2.04 0.395 2.68 0.485 ;
      LAYER MET2 ;
        RECT 2.45 0.625 2.55 1.16 ;
      LAYER VIA1 ;
        RECT 2.455 0.855 2.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.893 0.45 0.983 ;
      RECT 0.045 0.41 0.135 0.983 ;
      RECT 1.84 0.625 2.5 0.715 ;
      RECT 1.84 0.41 1.93 0.715 ;
      RECT 0.045 0.41 1.93 0.5 ;
      RECT 1.565 0.32 1.655 0.5 ;
      RECT 0.835 0.32 0.925 0.5 ;
      RECT 0.335 0.32 0.425 0.5 ;
      RECT 1.54 0.888 1.68 0.995 ;
      RECT 0.81 0.888 0.95 0.983 ;
      RECT 0.81 0.888 1.68 0.978 ;
      RECT 0.06 1.073 1.2 1.163 ;
      RECT 1.06 1.068 1.2 1.163 ;
  END
END OR3X8H7R

MACRO OR4X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X0P5H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.14 1.08 1.28 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.135 -0.08 1.275 0.175 ;
        RECT 0.57 -0.08 0.71 0.175 ;
        RECT 0.07 -0.08 0.16 0.375 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.995 0.6 1.145 0.78 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.625 0.79 0.775 ;
        RECT 0.7 0.55 0.79 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.41 0.455 0.59 0.545 ;
        RECT 0.41 0.455 0.56 0.63 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.435 0.24 1.545 1.08 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.895 0.185 1.085 ;
      RECT 0.045 0.895 1.345 0.985 ;
      RECT 1.255 0.265 1.345 0.985 ;
      RECT 0.295 0.265 1.345 0.355 ;
  END
END OR4X0P5H7R

MACRO OR4X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X0P7H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.14 1.09 1.28 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.135 -0.08 1.275 0.34 ;
        RECT 0.57 -0.08 0.71 0.34 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.625 1.145 0.78 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.625 0.835 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.36 0.625 0.56 0.79 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.435 0.249 1.545 1.145 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.91 0.185 1.12 ;
      RECT 0.045 0.91 1.345 1 ;
      RECT 1.255 0.445 1.345 1 ;
      RECT 0.295 0.445 1.345 0.535 ;
      RECT 0.86 0.265 1 0.535 ;
      RECT 0.295 0.265 0.435 0.535 ;
  END
END OR4X0P7H7R

MACRO OR4X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X1H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.115 1.06 1.255 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.125 -0.08 1.275 0.185 ;
        RECT 0.555 -0.08 0.705 0.185 ;
        RECT 0.07 -0.08 0.16 0.39 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.625 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.7 0.455 0.794 0.675 ;
        RECT 0.625 0.455 0.794 0.545 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.38 0.625 0.56 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.43 0.31 1.545 1.115 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.88 0.16 1.08 ;
      RECT 0.07 0.88 1.34 0.97 ;
      RECT 1.25 0.275 1.34 0.97 ;
      RECT 0.295 0.275 1.34 0.365 ;
  END
END OR4X1H7R

MACRO OR4X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X1P4H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.075 1.077 1.215 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.085 -0.08 1.235 0.185 ;
        RECT 0.555 -0.08 0.705 0.185 ;
        RECT 0.07 -0.08 0.16 0.39 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.625 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.455 0.85 0.575 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.365 0.625 0.545 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.43 0.31 1.545 1.012 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.897 1.34 0.987 ;
      RECT 1.25 0.275 1.34 0.987 ;
      RECT 0.295 0.275 1.34 0.365 ;
  END
END OR4X1P4H7R

MACRO OR4X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X2H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.665 1.01 1.755 1.48 ;
        RECT 1.115 1.06 1.255 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.665 -0.08 1.755 0.415 ;
        RECT 1.14 -0.08 1.23 0.21 ;
        RECT 0.6 -0.08 0.69 0.21 ;
        RECT 0.07 -0.08 0.16 0.415 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.975 0.615 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.825 0.835 0.975 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.48 0.545 0.78 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.415 0.275 1.545 1.15 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.06 1.065 1.015 1.155 ;
      RECT 0.925 0.865 1.015 1.155 ;
      RECT 0.925 0.865 1.325 0.955 ;
      RECT 1.235 0.3 1.325 0.955 ;
      RECT 0.31 0.3 1.325 0.39 ;
  END
END OR4X2H7R

MACRO OR4X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X3H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.665 1.035 1.755 1.48 ;
        RECT 1.1 1.05 1.19 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.665 -0.08 1.755 0.37 ;
        RECT 1.115 -0.08 1.205 0.24 ;
        RECT 0.585 -0.08 0.675 0.24 ;
        RECT 0.07 -0.08 0.16 0.37 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.975 0.615 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.655 0.625 0.805 0.805 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.675 0.545 0.975 ;
      LAYER MET2 ;
        RECT 0.45 0.63 0.55 1.16 ;
      LAYER VIA1 ;
        RECT 0.455 0.855 0.545 0.945 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.415 0.32 1.545 1.025 ;
      LAYER MET2 ;
        RECT 1.45 0.63 1.55 1.16 ;
      LAYER VIA1 ;
        RECT 1.455 0.855 1.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 1.065 0.985 1.155 ;
      RECT 0.895 0.865 0.985 1.155 ;
      RECT 0.07 1.015 0.16 1.155 ;
      RECT 0.895 0.865 1.325 0.955 ;
      RECT 1.235 0.33 1.325 0.955 ;
      RECT 0.295 0.33 1.325 0.42 ;
  END
END OR4X3H7R

MACRO OR4X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X4H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 1.805 1.075 1.945 1.48 ;
        RECT 1.115 1.045 1.255 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 1.805 -0.08 1.945 0.325 ;
        RECT 1.29 -0.08 1.43 0.34 ;
        RECT 1.085 -0.08 1.175 0.345 ;
        RECT 0.585 -0.08 0.675 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.965 0.625 1.145 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.855 0.775 0.945 ;
        RECT 0.685 0.665 0.775 0.945 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.365 0.625 0.545 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.54 0.895 2.345 0.985 ;
        RECT 2.255 0.415 2.345 0.985 ;
        RECT 1.54 0.415 2.345 0.505 ;
        RECT 2.085 0.235 2.225 0.505 ;
        RECT 2.11 0.895 2.2 1.195 ;
        RECT 1.54 0.265 1.68 0.505 ;
      LAYER MET2 ;
        RECT 2.25 0.63 2.35 1.16 ;
      LAYER VIA1 ;
        RECT 2.255 0.855 2.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.06 1.035 1.025 1.125 ;
      RECT 0.935 0.865 1.025 1.125 ;
      RECT 0.935 0.865 1.325 0.955 ;
      RECT 1.235 0.445 1.325 0.955 ;
      RECT 1.235 0.595 1.995 0.685 ;
      RECT 0.335 0.445 1.325 0.535 ;
      RECT 0.835 0.32 0.925 0.535 ;
      RECT 0.335 0.32 0.425 0.535 ;
  END
END OR4X4H7R

MACRO OR4X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X6H7R 0 0 ;
  SIZE 2.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.8 1.48 ;
        RECT 2.46 1.035 2.6 1.48 ;
        RECT 1.93 1.08 2.07 1.48 ;
        RECT 1.375 1.08 1.515 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.8 0.08 ;
        RECT 2.596 -0.08 2.686 0.345 ;
        RECT 2.056 -0.08 2.196 0.345 ;
        RECT 1.566 -0.08 1.656 0.345 ;
        RECT 1.336 -0.08 1.426 0.345 ;
        RECT 0.836 -0.08 0.926 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.19 0.62 1.375 0.77 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.855 1.01 0.945 ;
        RECT 0.92 0.615 1.01 0.945 ;
      LAYER MET2 ;
        RECT 0.85 0.625 0.95 1.16 ;
      LAYER VIA1 ;
        RECT 0.855 0.855 0.945 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.62 0.615 0.8 0.765 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.22 0.615 0.51 0.755 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.791 0.435 2.461 0.525 ;
        RECT 2.321 0.32 2.461 0.525 ;
        RECT 2.205 0.885 2.345 1.11 ;
        RECT 2.255 0.435 2.345 1.11 ;
        RECT 1.665 0.885 2.345 0.975 ;
        RECT 1.791 0.32 1.931 0.525 ;
        RECT 1.665 0.885 1.805 1.105 ;
      LAYER MET2 ;
        RECT 2.25 0.63 2.35 1.16 ;
      LAYER VIA1 ;
        RECT 2.255 0.855 2.345 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 1.035 1.19 1.125 ;
      RECT 1.1 0.9 1.19 1.125 ;
      RECT 1.1 0.9 1.575 0.99 ;
      RECT 1.485 0.435 1.575 0.99 ;
      RECT 1.485 0.615 2.135 0.705 ;
      RECT 0.07 0.435 1.575 0.525 ;
      RECT 1.086 0.37 1.176 0.525 ;
      RECT 0.57 0.22 0.66 0.525 ;
      RECT 0.07 0.205 0.16 0.525 ;
  END
END OR4X6H7R

MACRO SDFFNQX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNQX1H7R 0 0 ;
  SIZE 6.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.8 1.48 ;
        RECT 6.21 1.005 6.3 1.48 ;
        RECT 5.245 1.1 5.385 1.48 ;
        RECT 3.625 1.24 3.765 1.48 ;
        RECT 2.68 1.22 2.82 1.48 ;
        RECT 1.21 1.18 1.3 1.48 ;
        RECT 0.07 1.03 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.8 0.08 ;
        RECT 6.255 -0.08 6.345 0.375 ;
        RECT 4.92 -0.08 5.06 0.165 ;
        RECT 3.615 -0.08 3.755 0.165 ;
        RECT 2.65 -0.08 2.79 0.165 ;
        RECT 1.045 -0.08 1.185 0.165 ;
        RECT 0.07 -0.08 0.16 0.37 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.305 0.645 3.575 0.745 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.425 1.055 6.615 1.145 ;
        RECT 6.525 0.245 6.615 1.145 ;
      LAYER MET2 ;
        RECT 6.45 0.84 6.55 1.22 ;
      LAYER VIA1 ;
        RECT 6.455 1.055 6.545 1.145 ;
    END
  END Q
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.64 1.42 0.73 ;
        RECT 1.33 0.59 1.42 0.73 ;
        RECT 0.625 0.455 0.775 0.73 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.875 0.455 1.175 0.545 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.94 0.23 6.03 1.145 ;
      RECT 5.01 0.695 6.03 0.785 ;
      RECT 4.34 0.78 4.525 0.87 ;
      RECT 4.34 0.255 4.43 0.87 ;
      RECT 5.7 0.17 5.84 0.605 ;
      RECT 4.34 0.255 5.295 0.345 ;
      RECT 5.2 0.17 5.84 0.26 ;
      RECT 3.86 1.14 4.92 1.23 ;
      RECT 4.83 0.49 4.92 1.23 ;
      RECT 2.285 1.04 2.375 1.225 ;
      RECT 5.65 0.92 5.74 1.145 ;
      RECT 3.86 1.04 3.95 1.23 ;
      RECT 1.925 1.04 3.95 1.13 ;
      RECT 1.925 0.435 2.015 1.13 ;
      RECT 4.83 0.92 5.74 1.01 ;
      RECT 4.52 0.49 5.595 0.58 ;
      RECT 5.455 0.35 5.595 0.58 ;
      RECT 4.04 0.96 4.74 1.05 ;
      RECT 4.65 0.72 4.74 1.05 ;
      RECT 4.04 0.86 4.13 1.05 ;
      RECT 3.31 0.86 4.13 0.95 ;
      RECT 3.945 0.255 4.035 0.95 ;
      RECT 2.285 0.255 2.375 0.58 ;
      RECT 3.945 0.465 4.135 0.555 ;
      RECT 3.325 0.255 4.035 0.345 ;
      RECT 2.285 0.255 2.985 0.345 ;
      RECT 2.895 0.17 3.465 0.26 ;
      RECT 3.055 0.46 3.195 0.95 ;
      RECT 2.53 0.46 3.855 0.55 ;
      RECT 3.08 0.35 3.22 0.55 ;
      RECT 2.105 0.86 2.965 0.95 ;
      RECT 2.875 0.68 2.965 0.95 ;
      RECT 2.105 0.255 2.195 0.95 ;
      RECT 2.045 0.255 2.195 0.345 ;
      RECT 1.745 0.18 1.835 1.225 ;
      RECT 0.525 1 1.835 1.09 ;
      RECT 1.745 0.18 1.905 0.345 ;
      RECT 0.535 0.255 1.425 0.345 ;
      RECT 1.335 0.18 1.905 0.27 ;
      RECT 0.42 0.82 1.655 0.91 ;
      RECT 1.515 0.36 1.655 0.91 ;
      RECT 0.42 0.45 0.51 0.91 ;
  END
END SDFFNQX1H7R

MACRO SDFFNQX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNQX2H7R 0 0 ;
  SIZE 7 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7 1.48 ;
        RECT 6.75 1.005 6.84 1.48 ;
        RECT 6.21 1.03 6.3 1.48 ;
        RECT 5.245 1.055 5.385 1.48 ;
        RECT 3.625 1.235 3.765 1.48 ;
        RECT 2.68 1.22 2.82 1.48 ;
        RECT 1.24 1.18 1.33 1.48 ;
        RECT 0.07 1.025 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7 0.08 ;
        RECT 6.75 -0.08 6.84 0.37 ;
        RECT 6.21 -0.08 6.3 0.355 ;
        RECT 4.92 -0.08 5.06 0.165 ;
        RECT 3.615 -0.08 3.755 0.165 ;
        RECT 2.65 -0.08 2.79 0.165 ;
        RECT 1.045 -0.08 1.185 0.165 ;
        RECT 0.07 -0.08 0.16 0.37 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.305 0.645 3.575 0.745 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.455 0.245 6.57 1.1 ;
      LAYER MET2 ;
        RECT 6.45 0.425 6.55 0.96 ;
      LAYER VIA1 ;
        RECT 6.455 0.655 6.545 0.745 ;
    END
  END Q
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.625 0.64 1.42 0.73 ;
        RECT 1.33 0.57 1.42 0.73 ;
        RECT 0.625 0.455 0.775 0.73 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.875 0.455 1.175 0.545 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.95 0.23 6.04 1.145 ;
      RECT 5.01 0.695 6.04 0.785 ;
      RECT 4.34 0.78 4.525 0.87 ;
      RECT 4.34 0.255 4.43 0.87 ;
      RECT 5.77 0.17 5.86 0.605 ;
      RECT 4.34 0.255 5.295 0.345 ;
      RECT 5.2 0.17 5.86 0.26 ;
      RECT 3.86 1.14 4.92 1.23 ;
      RECT 4.83 0.44 4.92 1.23 ;
      RECT 2.285 1.04 2.375 1.225 ;
      RECT 5.65 0.875 5.74 1.145 ;
      RECT 3.86 1.04 3.95 1.23 ;
      RECT 1.925 1.04 3.95 1.13 ;
      RECT 1.925 0.435 2.015 1.13 ;
      RECT 4.83 0.875 5.74 0.965 ;
      RECT 4.52 0.44 5.595 0.53 ;
      RECT 5.455 0.35 5.595 0.53 ;
      RECT 4.04 0.96 4.74 1.05 ;
      RECT 4.65 0.74 4.74 1.05 ;
      RECT 4.04 0.255 4.13 1.05 ;
      RECT 3.31 0.86 4.13 0.95 ;
      RECT 2.285 0.255 2.375 0.58 ;
      RECT 3.325 0.255 4.13 0.345 ;
      RECT 2.285 0.255 2.985 0.345 ;
      RECT 2.895 0.18 3.465 0.27 ;
      RECT 3.055 0.46 3.195 0.95 ;
      RECT 3.76 0.46 3.85 0.745 ;
      RECT 2.53 0.46 3.85 0.55 ;
      RECT 3.08 0.36 3.22 0.55 ;
      RECT 2.105 0.86 2.965 0.95 ;
      RECT 2.875 0.67 2.965 0.95 ;
      RECT 2.105 0.255 2.195 0.95 ;
      RECT 2.035 0.255 2.195 0.345 ;
      RECT 1.745 0.17 1.835 1.225 ;
      RECT 0.525 1 1.835 1.09 ;
      RECT 1.745 0.17 1.91 0.345 ;
      RECT 0.525 0.255 1.425 0.345 ;
      RECT 1.335 0.17 1.91 0.26 ;
      RECT 0.42 0.82 1.655 0.91 ;
      RECT 1.515 0.36 1.655 0.91 ;
      RECT 0.42 0.46 0.51 0.91 ;
  END
END SDFFNQX2H7R

MACRO SDFFNQX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNQX3H7R 0 0 ;
  SIZE 6.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.6 1.48 ;
        RECT 6.27 1.04 6.36 1.48 ;
        RECT 5.76 1.04 5.85 1.48 ;
        RECT 4.895 1.11 5.035 1.48 ;
        RECT 3.625 1.24 3.765 1.48 ;
        RECT 2.7 1.24 2.84 1.48 ;
        RECT 1.24 1.24 1.38 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.6 0.08 ;
        RECT 6.405 -0.08 6.495 0.37 ;
        RECT 5.905 -0.08 5.995 0.37 ;
        RECT 4.895 -0.08 5.035 0.16 ;
        RECT 3.66 -0.08 3.75 0.2 ;
        RECT 2.69 -0.08 2.83 0.16 ;
        RECT 1.14 -0.08 1.28 0.16 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.38 0.65 3.605 0.77 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.26 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.02 0.655 6.245 0.745 ;
        RECT 6.155 0.29 6.245 0.745 ;
        RECT 6.02 0.655 6.11 1.05 ;
      LAYER MET2 ;
        RECT 6.05 0.43 6.15 0.96 ;
      LAYER VIA1 ;
        RECT 6.055 0.655 6.145 0.745 ;
    END
  END Q
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.365 0.445 1.455 0.755 ;
        RECT 0.655 0.445 1.455 0.535 ;
        RECT 0.655 0.425 0.81 0.605 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.625 1.235 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.49 0.69 5.58 1.095 ;
      RECT 5.49 0.69 5.745 0.785 ;
      RECT 5.655 0.295 5.745 0.785 ;
      RECT 4.745 0.69 5.745 0.78 ;
      RECT 4.325 0.255 4.415 0.99 ;
      RECT 4.325 0.255 5.114 0.345 ;
      RECT 4.325 0.255 5.161 0.299 ;
      RECT 4.325 0.255 5.199 0.279 ;
      RECT 5.16 0.17 5.56 0.26 ;
      RECT 5.076 0.236 5.56 0.26 ;
      RECT 5.114 0.194 5.16 0.322 ;
      RECT 4.12 1.14 4.595 1.23 ;
      RECT 4.505 0.46 4.595 1.23 ;
      RECT 1.965 1.14 2.5 1.23 ;
      RECT 2.41 1.06 4.21 1.15 ;
      RECT 1.965 0.48 2.055 1.23 ;
      RECT 4.505 0.93 5.325 1.02 ;
      RECT 4.505 0.46 5.355 0.55 ;
      RECT 5.265 0.35 5.355 0.55 ;
      RECT 5.265 0.35 5.405 0.44 ;
      RECT 3.33 0.88 4.03 0.97 ;
      RECT 3.94 0.29 4.03 0.97 ;
      RECT 2.355 0.25 2.445 0.635 ;
      RECT 3.37 0.29 4.235 0.38 ;
      RECT 4.03 0.17 4.235 0.38 ;
      RECT 2.355 0.25 3.01 0.34 ;
      RECT 3.37 0.17 3.46 0.38 ;
      RECT 2.92 0.17 3.46 0.26 ;
      RECT 3.03 0.87 3.215 0.96 ;
      RECT 3.125 0.35 3.215 0.96 ;
      RECT 3.76 0.47 3.85 0.655 ;
      RECT 3.125 0.47 3.85 0.56 ;
      RECT 3.1 0.35 3.24 0.55 ;
      RECT 2.56 0.46 3.24 0.55 ;
      RECT 2.175 0.223 2.265 1.05 ;
      RECT 2.175 0.74 2.815 0.83 ;
      RECT 2.725 0.685 3.035 0.775 ;
      RECT 0.66 1.06 1.875 1.15 ;
      RECT 1.785 0.17 1.875 1.15 ;
      RECT 1.785 0.17 1.91 0.37 ;
      RECT 0.855 0.25 1.46 0.34 ;
      RECT 0.61 0.245 0.945 0.335 ;
      RECT 1.37 0.17 1.91 0.26 ;
      RECT 0.87 0.88 1.69 0.97 ;
      RECT 1.6 0.35 1.69 0.97 ;
      RECT 0.87 0.725 0.96 0.97 ;
      RECT 0.43 0.725 0.96 0.815 ;
      RECT 0.43 0.475 0.52 0.815 ;
      RECT 1.55 0.35 1.69 0.44 ;
  END
END SDFFNQX3H7R

MACRO SDFFNRX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNRX0P5H7R 0 0 ;
  SIZE 7.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7.6 1.48 ;
        RECT 7.01 1.055 7.1 1.48 ;
        RECT 6.51 1.07 6.6 1.48 ;
        RECT 5.445 1.24 5.585 1.48 ;
        RECT 2.935 1.24 3.075 1.48 ;
        RECT 1.49 1.175 1.63 1.48 ;
        RECT 0.34 1.07 0.43 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7.6 0.08 ;
        RECT 7.055 -0.08 7.145 0.365 ;
        RECT 6.555 -0.08 6.645 0.355 ;
        RECT 5.575 -0.08 5.665 0.285 ;
        RECT 5.025 -0.08 5.115 0.33 ;
        RECT 3.7 -0.08 3.79 0.35 ;
        RECT 2.935 -0.08 3.075 0.16 ;
        RECT 1.32 -0.08 1.46 0.185 ;
        RECT 0.34 -0.08 0.43 0.33 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.565 0.625 1.745 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.415 0.61 0.595 0.76 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.25 0.95 7.44 1.04 ;
        RECT 7.35 0.225 7.44 1.04 ;
        RECT 7.255 0.225 7.44 0.38 ;
      LAYER MET2 ;
        RECT 7.25 0.18 7.35 0.56 ;
      LAYER VIA1 ;
        RECT 7.255 0.255 7.345 0.345 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.15 0.35 6.285 0.49 ;
        RECT 6.055 0.825 6.24 1.04 ;
        RECT 6.15 0.35 6.24 1.04 ;
      LAYER MET2 ;
        RECT 6.05 0.63 6.15 1.16 ;
      LAYER VIA1 ;
        RECT 6.055 0.855 6.145 0.945 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.625 0.745 5.775 0.945 ;
      LAYER MET2 ;
        RECT 5.65 0.625 5.75 1.16 ;
      LAYER VIA1 ;
        RECT 5.655 0.855 5.745 0.945 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.855 0.805 0.945 ;
        RECT 0.715 0.74 0.805 0.945 ;
        RECT 0.225 0.71 0.315 0.945 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.19 0.455 1.28 0.605 ;
        RECT 1.025 0.455 1.28 0.545 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.675 1.13 6.42 1.22 ;
      RECT 6.33 0.89 6.42 1.22 ;
      RECT 5.385 1.06 5.765 1.15 ;
      RECT 6.78 0.34 6.87 1.065 ;
      RECT 5.385 0.825 5.475 1.15 ;
      RECT 6.33 0.89 6.87 0.98 ;
      RECT 5.024 0.825 5.475 0.915 ;
      RECT 6.78 0.66 7.26 0.75 ;
      RECT 7.17 0.61 7.26 0.75 ;
      RECT 6.78 0.34 6.94 0.43 ;
      RECT 4.665 0.91 4.755 1.05 ;
      RECT 4.665 0.91 4.92 1 ;
      RECT 4.83 0.215 4.92 1 ;
      RECT 6.375 0.575 6.515 0.665 ;
      RECT 6.375 0.17 6.465 0.665 ;
      RECT 4.83 0.42 5.28 0.51 ;
      RECT 5.755 0.17 5.845 0.475 ;
      RECT 5.19 0.385 5.845 0.475 ;
      RECT 5.33 0.29 5.42 0.475 ;
      RECT 4.52 0.215 4.92 0.305 ;
      RECT 5.755 0.17 6.465 0.26 ;
      RECT 5.875 0.565 5.965 1.04 ;
      RECT 5.355 0.565 5.445 0.71 ;
      RECT 5.355 0.565 6.04 0.655 ;
      RECT 5.95 0.35 6.04 0.655 ;
      RECT 3.57 1.14 5.24 1.23 ;
      RECT 5.15 1.05 5.24 1.23 ;
      RECT 3.57 1.09 3.66 1.23 ;
      RECT 3.771 0.96 4.34 1.05 ;
      RECT 4.25 0.85 4.34 1.05 ;
      RECT 3.729 0.901 3.771 1.029 ;
      RECT 3.691 0.96 4.34 0.989 ;
      RECT 2.47 0.88 3.729 0.97 ;
      RECT 2.47 0.941 3.809 0.97 ;
      RECT 4.25 0.85 4.482 0.94 ;
      RECT 4.25 0.85 4.541 0.904 ;
      RECT 2.47 0.665 2.56 0.97 ;
      RECT 4.495 0.445 4.585 0.859 ;
      RECT 4.444 0.831 4.585 0.859 ;
      RECT 4.482 0.805 4.495 0.934 ;
      RECT 2.47 0.665 2.82 0.755 ;
      RECT 2.73 0.43 2.82 0.755 ;
      RECT 4.495 0.445 4.74 0.535 ;
      RECT 4.65 0.395 4.74 0.535 ;
      RECT 2.73 0.43 3.43 0.52 ;
      RECT 3.34 0.38 3.43 0.52 ;
      RECT 3.855 0.67 3.995 0.87 ;
      RECT 2.91 0.67 4.405 0.76 ;
      RECT 4.315 0.255 4.405 0.76 ;
      RECT 2.91 0.62 3 0.76 ;
      RECT 3.925 0.255 4.405 0.345 ;
      RECT 1.835 0.493 1.925 0.92 ;
      RECT 1.835 0.565 1.995 0.705 ;
      RECT 4.135 0.44 4.225 0.58 ;
      RECT 2.55 0.17 2.64 0.555 ;
      RECT 3.52 0.44 4.225 0.53 ;
      RECT 1.815 0.17 1.915 0.526 ;
      RECT 3.52 0.17 3.61 0.53 ;
      RECT 1.65 0.255 1.915 0.345 ;
      RECT 2.55 0.25 3.255 0.34 ;
      RECT 3.165 0.17 3.61 0.26 ;
      RECT 1.815 0.17 2.64 0.26 ;
      RECT 3.37 1.06 3.46 1.225 ;
      RECT 2.275 1.06 3.46 1.15 ;
      RECT 2.275 0.36 2.365 1.15 ;
      RECT 2.275 0.36 2.455 0.45 ;
      RECT 1.752 1.08 2.185 1.17 ;
      RECT 2.095 0.36 2.185 1.17 ;
      RECT 1.706 1.018 1.752 1.146 ;
      RECT 1.668 1.08 2.185 1.104 ;
      RECT 0.9 0.995 1.706 1.085 ;
      RECT 0.9 1.061 1.791 1.085 ;
      RECT 0.9 1.041 1.753 1.085 ;
      RECT 1.37 0.275 1.46 1.085 ;
      RECT 2.005 0.36 2.185 0.45 ;
      RECT 1.08 0.275 1.46 0.365 ;
      RECT 0.8 0.235 1.17 0.325 ;
      RECT 0.045 1.035 0.16 1.175 ;
      RECT 0.045 0.255 0.135 1.175 ;
      RECT 1.036 0.75 1.27 0.84 ;
      RECT 1.02 0.704 1.036 0.832 ;
      RECT 0.974 0.673 1.02 0.801 ;
      RECT 0.928 0.627 0.974 0.755 ;
      RECT 0.928 0.731 1.074 0.755 ;
      RECT 0.882 0.581 0.928 0.709 ;
      RECT 0.836 0.535 0.882 0.663 ;
      RECT 0.715 0.489 0.836 0.64 ;
      RECT 0.706 0.489 0.836 0.515 ;
      RECT 0.045 0.42 0.744 0.51 ;
      RECT 0.045 0.443 0.79 0.51 ;
      RECT 0.045 0.255 0.16 0.51 ;
  END
END SDFFNRX0P5H7R

MACRO SDFFNRX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNRX1H7R 0 0 ;
  SIZE 7.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7.6 1.48 ;
        RECT 7.01 1.055 7.1 1.48 ;
        RECT 6.51 1.065 6.6 1.48 ;
        RECT 5.445 1.24 5.585 1.48 ;
        RECT 2.875 1.24 3.015 1.48 ;
        RECT 1.5 1.15 1.59 1.48 ;
        RECT 0.34 1.07 0.43 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7.6 0.08 ;
        RECT 7.055 -0.08 7.145 0.345 ;
        RECT 6.555 -0.08 6.645 0.355 ;
        RECT 5.575 -0.08 5.665 0.23 ;
        RECT 5.025 -0.08 5.115 0.33 ;
        RECT 3.755 -0.08 3.845 0.35 ;
        RECT 2.935 -0.08 3.075 0.16 ;
        RECT 1.32 -0.08 1.46 0.185 ;
        RECT 0.34 -0.08 0.43 0.33 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.565 0.625 1.745 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.405 0.615 0.585 0.765 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.25 0.89 7.44 0.98 ;
        RECT 7.35 0.225 7.44 0.98 ;
        RECT 7.255 0.225 7.44 0.375 ;
      LAYER MET2 ;
        RECT 7.25 0.18 7.35 0.56 ;
      LAYER VIA1 ;
        RECT 7.255 0.255 7.345 0.345 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.15 0.35 6.285 0.49 ;
        RECT 6.055 0.825 6.24 1.015 ;
        RECT 6.15 0.35 6.24 1.015 ;
      LAYER MET2 ;
        RECT 6.05 0.63 6.15 1.16 ;
      LAYER VIA1 ;
        RECT 6.055 0.855 6.145 0.945 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.625 0.745 5.775 0.945 ;
      LAYER MET2 ;
        RECT 5.65 0.625 5.75 1.16 ;
      LAYER VIA1 ;
        RECT 5.655 0.855 5.745 0.945 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.855 0.805 0.945 ;
        RECT 0.715 0.74 0.805 0.945 ;
        RECT 0.225 0.715 0.315 0.945 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.19 0.455 1.28 0.605 ;
        RECT 1.025 0.455 1.28 0.545 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.675 1.13 6.42 1.22 ;
      RECT 6.33 0.785 6.42 1.22 ;
      RECT 5.385 1.06 5.765 1.15 ;
      RECT 6.78 0.34 6.87 1.065 ;
      RECT 5.385 0.83 5.475 1.15 ;
      RECT 5.01 0.83 5.475 0.92 ;
      RECT 6.33 0.785 6.87 0.875 ;
      RECT 6.78 0.66 7.26 0.75 ;
      RECT 7.17 0.61 7.26 0.75 ;
      RECT 6.78 0.34 6.92 0.43 ;
      RECT 4.675 0.91 4.765 1.05 ;
      RECT 4.675 0.91 4.92 1 ;
      RECT 4.83 0.215 4.92 1 ;
      RECT 6.375 0.575 6.535 0.665 ;
      RECT 6.375 0.17 6.465 0.665 ;
      RECT 4.83 0.42 5.295 0.51 ;
      RECT 5.205 0.32 5.295 0.51 ;
      RECT 5.205 0.32 5.845 0.41 ;
      RECT 5.755 0.17 5.845 0.41 ;
      RECT 4.53 0.215 4.92 0.305 ;
      RECT 5.755 0.17 6.465 0.26 ;
      RECT 5.875 0.555 5.965 1.04 ;
      RECT 5.385 0.555 5.475 0.71 ;
      RECT 5.385 0.555 6.04 0.645 ;
      RECT 5.95 0.35 6.04 0.645 ;
      RECT 3.57 1.14 5.255 1.23 ;
      RECT 5.165 1.05 5.255 1.23 ;
      RECT 3.57 1.09 3.66 1.23 ;
      RECT 3.771 0.96 4.34 1.05 ;
      RECT 3.729 0.901 3.771 1.029 ;
      RECT 3.691 0.96 4.34 0.989 ;
      RECT 2.73 0.88 3.729 0.97 ;
      RECT 4.485 0.445 4.575 0.965 ;
      RECT 4.25 0.875 4.575 0.965 ;
      RECT 2.73 0.941 3.809 0.97 ;
      RECT 2.73 0.43 2.82 0.97 ;
      RECT 2.445 0.695 2.82 0.785 ;
      RECT 4.485 0.445 4.74 0.535 ;
      RECT 4.65 0.395 4.74 0.535 ;
      RECT 2.73 0.43 3.46 0.52 ;
      RECT 3.37 0.35 3.46 0.52 ;
      RECT 3.91 0.695 4.05 0.87 ;
      RECT 2.91 0.695 4.395 0.785 ;
      RECT 4.305 0.215 4.395 0.785 ;
      RECT 2.91 0.645 3 0.785 ;
      RECT 4.01 0.215 4.395 0.305 ;
      RECT 1.795 0.875 1.995 0.965 ;
      RECT 1.905 0.559 1.995 0.965 ;
      RECT 1.903 0.49 1.905 0.618 ;
      RECT 4.125 0.44 4.215 0.6 ;
      RECT 1.857 0.466 1.903 0.594 ;
      RECT 1.857 0.514 1.951 0.594 ;
      RECT 2.55 0.17 2.64 0.555 ;
      RECT 1.811 0.42 1.857 0.548 ;
      RECT 3.575 0.44 4.215 0.53 ;
      RECT 1.765 0.374 1.811 0.502 ;
      RECT 1.721 0.17 1.765 0.457 ;
      RECT 3.575 0.17 3.665 0.53 ;
      RECT 1.675 0.17 1.765 0.412 ;
      RECT 2.55 0.25 3.255 0.34 ;
      RECT 3.165 0.17 3.665 0.26 ;
      RECT 1.675 0.17 2.64 0.26 ;
      RECT 3.37 1.06 3.46 1.225 ;
      RECT 2.265 1.06 3.46 1.15 ;
      RECT 2.265 0.36 2.355 1.15 ;
      RECT 2.265 0.36 2.455 0.45 ;
      RECT 1.715 1.055 2.175 1.145 ;
      RECT 2.085 0.36 2.175 1.145 ;
      RECT 1.669 0.993 1.715 1.121 ;
      RECT 1.631 1.055 2.175 1.079 ;
      RECT 0.98 0.97 1.669 1.06 ;
      RECT 0.98 1.036 1.754 1.06 ;
      RECT 0.98 1.016 1.716 1.06 ;
      RECT 1.37 0.275 1.46 1.06 ;
      RECT 2.005 0.36 2.175 0.45 ;
      RECT 1.08 0.275 1.46 0.365 ;
      RECT 0.8 0.26 1.17 0.35 ;
      RECT 0.045 1.03 0.185 1.12 ;
      RECT 0.045 0.255 0.135 1.12 ;
      RECT 1.041 0.75 1.27 0.84 ;
      RECT 1.025 0.704 1.041 0.832 ;
      RECT 0.979 0.673 1.025 0.801 ;
      RECT 0.933 0.627 0.979 0.755 ;
      RECT 0.933 0.731 1.079 0.755 ;
      RECT 0.887 0.581 0.933 0.709 ;
      RECT 0.841 0.535 0.887 0.663 ;
      RECT 0.69 0.496 0.841 0.64 ;
      RECT 0.045 0.435 0.764 0.525 ;
      RECT 0.045 0.458 0.81 0.525 ;
      RECT 0.045 0.255 0.16 0.525 ;
  END
END SDFFNRX1H7R

MACRO SDFFNRX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNRX2H7R 0 0 ;
  SIZE 7.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7.6 1.48 ;
        RECT 7.01 1.055 7.1 1.48 ;
        RECT 6.47 1.095 6.61 1.48 ;
        RECT 5.37 1.195 5.46 1.48 ;
        RECT 2.875 1.24 3.015 1.48 ;
        RECT 1.475 1.125 1.615 1.48 ;
        RECT 0.34 1.07 0.43 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7.6 0.08 ;
        RECT 7.005 -0.08 7.095 0.345 ;
        RECT 6.525 -0.08 6.615 0.33 ;
        RECT 5.545 -0.08 5.635 0.33 ;
        RECT 5.065 -0.08 5.155 0.33 ;
        RECT 3.685 -0.08 3.775 0.345 ;
        RECT 2.915 -0.08 3.055 0.16 ;
        RECT 1.32 -0.08 1.46 0.185 ;
        RECT 0.34 -0.08 0.43 0.33 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.565 0.625 1.745 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.405 0.615 0.585 0.765 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.25 0.83 7.395 0.92 ;
        RECT 7.305 0.225 7.395 0.92 ;
        RECT 7.255 0.225 7.395 0.375 ;
      LAYER MET2 ;
        RECT 7.25 0.18 7.35 0.56 ;
      LAYER VIA1 ;
        RECT 7.255 0.255 7.345 0.345 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.165 0.35 6.255 0.706 ;
        RECT 6.101 0.688 6.211 0.751 ;
        RECT 6.145 0.656 6.165 0.784 ;
        RECT 6.055 0.733 6.145 0.975 ;
      LAYER MET2 ;
        RECT 6.05 0.63 6.15 1.16 ;
      LAYER VIA1 ;
        RECT 6.055 0.855 6.145 0.945 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.575 0.61 5.775 0.745 ;
      LAYER MET2 ;
        RECT 5.65 0.425 5.75 0.96 ;
      LAYER VIA1 ;
        RECT 5.655 0.655 5.745 0.745 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.855 0.805 0.945 ;
        RECT 0.715 0.74 0.805 0.945 ;
        RECT 0.225 0.71 0.315 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.19 0.455 1.28 0.605 ;
        RECT 1.025 0.455 1.28 0.545 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.57 1.13 6.38 1.22 ;
      RECT 6.29 0.91 6.38 1.22 ;
      RECT 5.57 1.015 5.66 1.22 ;
      RECT 5.21 1.015 5.66 1.105 ;
      RECT 5.21 0.85 5.3 1.105 ;
      RECT 6.29 0.91 6.865 1 ;
      RECT 6.775 0.315 6.865 1 ;
      RECT 4.87 0.85 5.3 0.94 ;
      RECT 6.775 0.605 7.205 0.695 ;
      RECT 4.525 0.91 4.615 1.05 ;
      RECT 4.525 0.91 4.73 1 ;
      RECT 4.64 0.645 4.73 1 ;
      RECT 4.64 0.645 4.975 0.735 ;
      RECT 4.885 0.235 4.975 0.735 ;
      RECT 6.345 0.17 6.435 0.69 ;
      RECT 4.885 0.435 5.435 0.525 ;
      RECT 5.725 0.17 5.815 0.52 ;
      RECT 5.315 0.43 5.815 0.52 ;
      RECT 5.315 0.315 5.405 0.525 ;
      RECT 4.53 0.235 4.975 0.325 ;
      RECT 5.725 0.17 6.435 0.26 ;
      RECT 5.75 0.835 5.84 1.04 ;
      RECT 5.395 0.835 5.965 0.925 ;
      RECT 5.875 0.661 5.965 0.925 ;
      RECT 5.395 0.62 5.485 0.925 ;
      RECT 5.165 0.62 5.485 0.71 ;
      RECT 5.905 0.35 5.995 0.699 ;
      RECT 3.57 1.14 5.12 1.23 ;
      RECT 5.03 1.035 5.12 1.23 ;
      RECT 3.57 1.09 3.66 1.23 ;
      RECT 3.771 0.96 4.415 1.05 ;
      RECT 4.325 0.72 4.415 1.05 ;
      RECT 3.729 0.901 3.771 1.029 ;
      RECT 3.691 0.96 4.415 0.989 ;
      RECT 2.73 0.88 3.729 0.97 ;
      RECT 2.73 0.941 3.809 0.97 ;
      RECT 2.73 0.43 2.82 0.97 ;
      RECT 2.455 0.76 2.82 0.85 ;
      RECT 4.325 0.72 4.55 0.81 ;
      RECT 4.46 0.465 4.55 0.81 ;
      RECT 4.46 0.465 4.795 0.555 ;
      RECT 4.705 0.415 4.795 0.555 ;
      RECT 2.73 0.43 3.415 0.52 ;
      RECT 3.325 0.35 3.415 0.52 ;
      RECT 1.835 0.535 1.925 0.955 ;
      RECT 1.835 0.535 1.975 0.675 ;
      RECT 4.28 0.17 4.37 0.62 ;
      RECT 1.825 0.17 1.915 0.58 ;
      RECT 2.55 0.17 2.64 0.555 ;
      RECT 3.505 0.435 3.955 0.525 ;
      RECT 3.865 0.17 3.955 0.525 ;
      RECT 3.505 0.17 3.595 0.525 ;
      RECT 1.65 0.255 1.915 0.345 ;
      RECT 2.55 0.25 3.235 0.34 ;
      RECT 3.865 0.17 4.37 0.26 ;
      RECT 3.145 0.17 3.595 0.26 ;
      RECT 1.825 0.17 2.64 0.26 ;
      RECT 3.91 0.695 4.05 0.87 ;
      RECT 2.91 0.695 4.135 0.785 ;
      RECT 4.045 0.35 4.135 0.785 ;
      RECT 2.91 0.645 3 0.785 ;
      RECT 4.045 0.35 4.185 0.44 ;
      RECT 3.37 1.06 3.46 1.225 ;
      RECT 2.275 1.06 3.46 1.15 ;
      RECT 2.275 0.36 2.365 1.15 ;
      RECT 2.275 0.36 2.455 0.45 ;
      RECT 1.756 1.045 2.185 1.135 ;
      RECT 2.095 0.36 2.185 1.135 ;
      RECT 1.74 0.999 1.756 1.127 ;
      RECT 1.694 0.968 1.74 1.096 ;
      RECT 1.656 1.026 1.794 1.054 ;
      RECT 0.98 0.945 1.694 1.035 ;
      RECT 1.37 0.275 1.46 1.035 ;
      RECT 2.005 0.36 2.185 0.45 ;
      RECT 1.08 0.275 1.46 0.365 ;
      RECT 0.805 0.26 1.17 0.35 ;
      RECT 0.045 1.01 0.16 1.15 ;
      RECT 0.045 0.23 0.135 1.15 ;
      RECT 1.036 0.75 1.27 0.84 ;
      RECT 1.02 0.704 1.036 0.832 ;
      RECT 0.974 0.673 1.02 0.801 ;
      RECT 0.928 0.627 0.974 0.755 ;
      RECT 0.928 0.731 1.074 0.755 ;
      RECT 0.882 0.581 0.928 0.709 ;
      RECT 0.836 0.535 0.882 0.663 ;
      RECT 0.715 0.489 0.836 0.64 ;
      RECT 0.706 0.489 0.836 0.515 ;
      RECT 0.045 0.42 0.744 0.51 ;
      RECT 0.045 0.443 0.79 0.51 ;
      RECT 0.045 0.23 0.16 0.51 ;
  END
END SDFFNRX2H7R

MACRO SDFFNRX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNRX3H7R 0 0 ;
  SIZE 8.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 8.4 1.48 ;
        RECT 8.185 1.055 8.275 1.48 ;
        RECT 7.675 1.055 7.765 1.48 ;
        RECT 6.81 1.24 6.955 1.48 ;
        RECT 5.775 1.225 5.915 1.48 ;
        RECT 2.985 1.24 3.125 1.48 ;
        RECT 1.6 1.225 1.74 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 8.4 0.08 ;
        RECT 8.185 -0.08 8.275 0.345 ;
        RECT 7.675 -0.08 7.765 0.345 ;
        RECT 6.945 -0.08 7.035 0.355 ;
        RECT 5.965 -0.08 6.055 0.285 ;
        RECT 5.455 -0.08 5.545 0.345 ;
        RECT 3.895 -0.08 3.985 0.345 ;
        RECT 3.05 -0.08 3.19 0.16 ;
        RECT 1.465 -0.08 1.605 0.185 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.74 0.625 1.945 0.775 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.405 0.655 0.64 0.77 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.935 0.225 8.025 1.03 ;
        RECT 7.855 0.225 8.025 0.375 ;
      LAYER MET2 ;
        RECT 7.85 0.18 7.95 0.56 ;
      LAYER VIA1 ;
        RECT 7.855 0.255 7.945 0.345 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.195 0.25 7.285 1.045 ;
        RECT 6.505 0.855 7.285 0.945 ;
        RECT 6.585 0.35 6.675 0.945 ;
        RECT 6.505 0.855 6.595 1.045 ;
      LAYER MET2 ;
        RECT 6.65 0.625 6.75 1.16 ;
      LAYER VIA1 ;
        RECT 6.655 0.855 6.745 0.945 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.05 0.585 6.195 0.775 ;
      LAYER MET2 ;
        RECT 6.05 0.43 6.15 0.96 ;
      LAYER VIA1 ;
        RECT 6.055 0.655 6.145 0.745 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.865 0.995 0.955 ;
        RECT 0.905 0.735 0.995 0.955 ;
        RECT 0.225 0.855 0.375 0.955 ;
        RECT 0.225 0.65 0.315 0.955 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.26 0.455 1.425 0.585 ;
        RECT 1.205 0.455 1.425 0.56 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 6.005 1.14 6.674 1.23 ;
      RECT 7.069 1.135 7.515 1.225 ;
      RECT 7.425 0.315 7.515 1.225 ;
      RECT 7.032 1.078 7.069 1.207 ;
      RECT 6.994 1.135 7.515 1.169 ;
      RECT 6.005 1.14 6.754 1.169 ;
      RECT 6.716 1.06 7.032 1.15 ;
      RECT 6.674 1.081 6.716 1.209 ;
      RECT 6.005 1.045 6.095 1.23 ;
      RECT 5.69 1.045 6.095 1.135 ;
      RECT 6.636 1.121 7.107 1.15 ;
      RECT 7.069 1.116 7.107 1.225 ;
      RECT 5.69 0.87 5.78 1.135 ;
      RECT 5.34 0.87 5.43 1.01 ;
      RECT 5.34 0.87 5.78 0.96 ;
      RECT 7.425 0.66 7.845 0.75 ;
      RECT 7.755 0.61 7.845 0.75 ;
      RECT 4.63 0.91 4.72 1.05 ;
      RECT 4.63 0.91 5.082 1 ;
      RECT 4.63 0.91 5.128 0.977 ;
      RECT 5.044 0.891 5.174 0.931 ;
      RECT 5.082 0.849 5.174 0.931 ;
      RECT 5.082 0.849 5.22 0.885 ;
      RECT 5.128 0.803 5.225 0.86 ;
      RECT 5.174 0.757 5.271 0.834 ;
      RECT 5.22 0.731 5.225 0.86 ;
      RECT 5.225 0.23 5.315 0.789 ;
      RECT 6.765 0.575 6.95 0.665 ;
      RECT 6.765 0.17 6.855 0.665 ;
      RECT 5.225 0.435 5.825 0.525 ;
      RECT 5.735 0.23 5.825 0.525 ;
      RECT 6.145 0.17 6.235 0.465 ;
      RECT 5.735 0.375 6.235 0.465 ;
      RECT 4.95 0.23 5.315 0.32 ;
      RECT 6.145 0.17 6.855 0.26 ;
      RECT 6.185 0.865 6.275 1.04 ;
      RECT 5.87 0.865 6.415 0.955 ;
      RECT 6.325 0.35 6.415 0.955 ;
      RECT 5.87 0.62 5.96 0.955 ;
      RECT 5.61 0.62 5.96 0.71 ;
      RECT 3.725 1.14 5.6 1.23 ;
      RECT 5.46 1.095 5.6 1.23 ;
      RECT 3.725 1.07 3.815 1.23 ;
      RECT 3.923 0.96 4.54 1.05 ;
      RECT 4.45 0.73 4.54 1.05 ;
      RECT 3.881 0.901 3.923 1.029 ;
      RECT 3.843 0.96 4.54 0.989 ;
      RECT 2.6 0.88 3.881 0.97 ;
      RECT 2.6 0.941 3.961 0.97 ;
      RECT 2.795 0.635 2.885 0.97 ;
      RECT 2.6 0.815 2.69 0.97 ;
      RECT 4.45 0.73 5.006 0.82 ;
      RECT 4.968 0.711 5.091 0.758 ;
      RECT 5.006 0.672 5.045 0.801 ;
      RECT 5.045 0.41 5.135 0.713 ;
      RECT 2.795 0.635 2.931 0.673 ;
      RECT 2.865 0.43 2.955 0.638 ;
      RECT 2.841 0.6 2.955 0.638 ;
      RECT 2.865 0.43 3.58 0.52 ;
      RECT 3.49 0.35 3.58 0.52 ;
      RECT 1.865 0.87 2.15 0.96 ;
      RECT 2.06 0.536 2.15 0.96 ;
      RECT 4.69 0.55 4.86 0.64 ;
      RECT 4.77 0.17 4.86 0.64 ;
      RECT 3.695 0.49 4.175 0.58 ;
      RECT 4.085 0.17 4.175 0.58 ;
      RECT 2.016 0.446 2.06 0.574 ;
      RECT 2.685 0.17 2.775 0.55 ;
      RECT 2.016 0.491 2.106 0.574 ;
      RECT 1.97 0.401 2.016 0.529 ;
      RECT 3.695 0.17 3.785 0.58 ;
      RECT 1.926 0.17 1.97 0.484 ;
      RECT 1.88 0.17 1.97 0.439 ;
      RECT 2.685 0.25 3.4 0.34 ;
      RECT 4.085 0.17 4.86 0.26 ;
      RECT 3.31 0.17 3.785 0.26 ;
      RECT 1.88 0.17 2.775 0.26 ;
      RECT 3.999 0.7 4.139 0.87 ;
      RECT 3.01 0.7 4.244 0.79 ;
      RECT 3.01 0.7 4.29 0.767 ;
      RECT 4.206 0.681 4.356 0.701 ;
      RECT 4.29 0.606 4.31 0.734 ;
      RECT 4.244 0.639 4.356 0.701 ;
      RECT 4.31 0.35 4.4 0.656 ;
      RECT 4.31 0.35 4.64 0.44 ;
      RECT 3.525 1.06 3.615 1.225 ;
      RECT 2.42 1.06 3.615 1.15 ;
      RECT 2.42 0.35 2.51 1.15 ;
      RECT 2.42 0.35 2.59 0.44 ;
      RECT 1.836 1.095 2.33 1.185 ;
      RECT 2.24 0.35 2.33 1.185 ;
      RECT 1.824 1.051 1.836 1.179 ;
      RECT 1.786 1.095 2.33 1.154 ;
      RECT 1.105 1.045 1.824 1.135 ;
      RECT 1.105 1.076 1.874 1.135 ;
      RECT 1.515 0.275 1.605 1.135 ;
      RECT 2.17 0.35 2.33 0.44 ;
      RECT 0.925 0.275 1.605 0.365 ;
      RECT 0.045 1.075 0.185 1.165 ;
      RECT 0.045 0.295 0.135 1.165 ;
      RECT 1.1 0.75 1.395 0.84 ;
      RECT 1.1 0.651 1.19 0.84 ;
      RECT 1.072 0.569 1.1 0.697 ;
      RECT 1.034 0.606 1.146 0.664 ;
      RECT 0.87 0.555 1.072 0.645 ;
      RECT 0.87 0.455 0.96 0.645 ;
      RECT 0.045 0.455 0.96 0.545 ;
      RECT 0.045 0.295 0.16 0.545 ;
  END
END SDFFNRX3H7R

MACRO SDFFNSRX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNSRX0P5H7R 0 0 ;
  SIZE 8.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 8.4 1.48 ;
        RECT 7.915 0.855 8.005 1.48 ;
        RECT 7.145 1.095 7.285 1.48 ;
        RECT 6.316 1.225 6.456 1.48 ;
        RECT 5.305 1.225 5.445 1.48 ;
        RECT 2.835 1.24 2.975 1.48 ;
        RECT 1.505 1.24 1.645 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 8.4 0.08 ;
        RECT 7.56 -0.08 7.65 0.365 ;
        RECT 6.855 -0.08 6.995 0.26 ;
        RECT 5.95 -0.08 6.09 0.16 ;
        RECT 2.865 -0.08 3.005 0.16 ;
        RECT 1.395 -0.08 1.535 0.175 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.535 0.625 1.75 0.805 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.43 0.645 0.625 0.781 ;
        RECT 0.444 0.645 0.58 0.825 ;
        RECT 0.43 0.645 0.58 0.782 ;
        RECT 0.405 0.645 0.625 0.75 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 8.165 0.25 8.255 1.085 ;
        RECT 7.785 0.25 8.255 0.35 ;
      LAYER MET2 ;
        RECT 7.85 0.18 7.95 0.56 ;
      LAYER VIA1 ;
        RECT 7.855 0.255 7.945 0.345 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.555 0.645 7.645 1.05 ;
        RECT 7.38 0.645 7.645 0.735 ;
        RECT 7.38 0.25 7.47 0.735 ;
        RECT 7.17 0.25 7.47 0.35 ;
      LAYER MET2 ;
        RECT 7.25 0.18 7.35 0.56 ;
      LAYER VIA1 ;
        RECT 7.255 0.255 7.345 0.345 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.985 0.45 6.175 0.69 ;
      LAYER MET2 ;
        RECT 6.05 0.23 6.15 0.76 ;
      LAYER VIA1 ;
        RECT 6.055 0.455 6.145 0.545 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.715 0.74 0.805 0.906 ;
        RECT 0.646 0.896 0.761 0.951 ;
        RECT 0.684 0.861 0.715 0.99 ;
        RECT 0.281 0.915 0.684 1.005 ;
        RECT 0.225 0.825 0.35 0.972 ;
        RECT 0.225 0.715 0.315 0.972 ;
        RECT 0.271 0.915 0.684 1 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.435 1.265 0.565 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END SI
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.28 0.53 6.62 0.75 ;
      LAYER MET2 ;
        RECT 6.45 0.425 6.55 0.96 ;
      LAYER VIA1 ;
        RECT 6.455 0.655 6.545 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 7.375 1.14 7.825 1.23 ;
      RECT 7.735 0.62 7.825 1.23 ;
      RECT 6.589 1.14 7.01 1.23 ;
      RECT 6.92 0.915 7.01 1.23 ;
      RECT 5.58 1.14 6.183 1.23 ;
      RECT 6.578 1.096 6.589 1.225 ;
      RECT 5.569 1.096 5.58 1.225 ;
      RECT 4.88 1.07 4.97 1.225 ;
      RECT 6.532 1.068 6.578 1.196 ;
      RECT 5.523 1.068 5.569 1.196 ;
      RECT 4.88 1.07 5.239 1.16 ;
      RECT 4.88 1.07 5.264 1.148 ;
      RECT 7.375 0.915 7.465 1.23 ;
      RECT 6.494 1.121 6.627 1.154 ;
      RECT 6.145 1.121 6.278 1.154 ;
      RECT 6.229 1.05 6.24 1.179 ;
      RECT 5.485 1.121 5.618 1.154 ;
      RECT 6.24 1.045 6.532 1.135 ;
      RECT 5.226 1.045 5.523 1.135 ;
      RECT 6.183 1.079 6.229 1.207 ;
      RECT 5.201 1.057 5.239 1.16 ;
      RECT 6.92 0.915 7.465 1.005 ;
      RECT 7.2 0.44 7.29 1.005 ;
      RECT 7.735 0.62 8.075 0.71 ;
      RECT 6.75 0.44 7.29 0.53 ;
      RECT 6.605 0.35 6.84 0.44 ;
      RECT 6.605 0.205 6.695 0.44 ;
      RECT 6.665 0.865 6.83 1.05 ;
      RECT 6.74 0.62 6.83 1.05 ;
      RECT 5.656 0.96 6.107 1.05 ;
      RECT 4.52 0.71 4.61 1.05 ;
      RECT 5.645 0.916 5.656 1.045 ;
      RECT 5.645 0.96 6.153 1.027 ;
      RECT 5.599 0.888 5.645 1.016 ;
      RECT 6.069 0.941 6.202 0.974 ;
      RECT 6.153 0.87 6.164 0.999 ;
      RECT 5.561 0.941 5.694 0.974 ;
      RECT 6.164 0.865 6.83 0.955 ;
      RECT 5.2 0.865 5.599 0.955 ;
      RECT 6.107 0.899 6.83 0.955 ;
      RECT 5.2 0.71 5.29 0.955 ;
      RECT 4.52 0.71 5.29 0.8 ;
      RECT 6.74 0.62 7.11 0.71 ;
      RECT 4.915 0.35 5.005 0.8 ;
      RECT 4.38 0.35 5.495 0.44 ;
      RECT 3.595 0.17 3.685 0.381 ;
      RECT 5.873 0.25 6.49 0.34 ;
      RECT 5.831 0.191 5.873 0.319 ;
      RECT 5.793 0.25 6.49 0.279 ;
      RECT 3.595 0.17 5.831 0.26 ;
      RECT 3.595 0.231 5.911 0.26 ;
      RECT 5.805 0.78 6.03 0.87 ;
      RECT 5.805 0.53 5.895 0.87 ;
      RECT 5.155 0.53 5.895 0.62 ;
      RECT 5.615 0.35 5.755 0.62 ;
      RECT 3.48 1.14 4.79 1.23 ;
      RECT 4.7 0.89 4.79 1.23 ;
      RECT 3.48 1.07 3.57 1.23 ;
      RECT 4.7 0.89 5.11 0.98 ;
      RECT 3.678 0.96 4.43 1.05 ;
      RECT 4.34 0.53 4.43 1.05 ;
      RECT 3.636 0.901 3.678 1.029 ;
      RECT 3.598 0.96 4.43 0.989 ;
      RECT 2.5 0.88 3.636 0.97 ;
      RECT 2.5 0.941 3.716 0.97 ;
      RECT 2.5 0.43 2.59 0.97 ;
      RECT 4.34 0.53 4.825 0.62 ;
      RECT 2.5 0.43 3.295 0.52 ;
      RECT 3.205 0.35 3.295 0.52 ;
      RECT 3.754 0.78 4.25 0.87 ;
      RECT 4.16 0.35 4.25 0.87 ;
      RECT 3.712 0.721 3.754 0.849 ;
      RECT 3.674 0.78 4.25 0.809 ;
      RECT 2.705 0.7 3.712 0.79 ;
      RECT 2.705 0.761 3.792 0.79 ;
      RECT 3.985 0.35 4.25 0.44 ;
      RECT 1.785 0.905 1.95 0.995 ;
      RECT 1.86 0.535 1.95 0.995 ;
      RECT 3.821 0.58 4.07 0.67 ;
      RECT 3.799 0.531 3.821 0.659 ;
      RECT 3.761 0.58 4.07 0.629 ;
      RECT 3.39 0.52 3.799 0.61 ;
      RECT 3.39 0.561 3.859 0.61 ;
      RECT 1.821 0.446 1.86 0.575 ;
      RECT 1.821 0.523 1.929 0.575 ;
      RECT 1.775 0.404 1.821 0.532 ;
      RECT 1.775 0.489 1.906 0.532 ;
      RECT 3.39 0.17 3.48 0.61 ;
      RECT 1.731 0.17 1.775 0.487 ;
      RECT 1.685 0.17 1.775 0.442 ;
      RECT 2.685 0.25 3.081 0.34 ;
      RECT 2.685 0.25 3.161 0.279 ;
      RECT 3.123 0.17 3.48 0.26 ;
      RECT 3.043 0.231 3.48 0.26 ;
      RECT 3.081 0.191 3.123 0.319 ;
      RECT 1.685 0.17 2.775 0.26 ;
      RECT 3.27 1.06 3.36 1.225 ;
      RECT 2.29 1.06 3.36 1.15 ;
      RECT 2.29 0.35 2.38 1.15 ;
      RECT 2.225 0.35 2.38 0.44 ;
      RECT 1.763 1.14 2.13 1.23 ;
      RECT 2.04 0.35 2.13 1.23 ;
      RECT 1.721 1.081 1.763 1.209 ;
      RECT 1.683 1.14 2.13 1.169 ;
      RECT 0.76 1.06 1.721 1.15 ;
      RECT 0.76 1.121 1.801 1.15 ;
      RECT 1.355 0.335 1.445 1.15 ;
      RECT 1.975 0.35 2.13 0.44 ;
      RECT 1.349 0.264 1.355 0.392 ;
      RECT 1.303 0.238 1.349 0.366 ;
      RECT 1.303 0.29 1.401 0.366 ;
      RECT 1.265 0.29 1.401 0.324 ;
      RECT 0.755 0.215 1.303 0.305 ;
      RECT 0.045 1.08 0.185 1.17 ;
      RECT 0.045 0.395 0.135 1.17 ;
      RECT 1.028 0.735 1.235 0.825 ;
      RECT 1.026 0.696 1.028 0.824 ;
      RECT 0.98 0.672 1.026 0.8 ;
      RECT 0.934 0.626 0.98 0.754 ;
      RECT 0.934 0.716 1.066 0.754 ;
      RECT 0.888 0.58 0.934 0.708 ;
      RECT 0.842 0.534 0.888 0.662 ;
      RECT 0.796 0.488 0.842 0.616 ;
      RECT 0.758 0.534 0.888 0.574 ;
      RECT 0.445 0.465 0.796 0.555 ;
      RECT 0.045 0.395 0.535 0.485 ;
      RECT 0.07 0.224 0.16 0.485 ;
  END
END SDFFNSRX0P5H7R

MACRO SDFFNSRX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNSRX1H7R 0 0 ;
  SIZE 8.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 8.4 1.48 ;
        RECT 7.915 0.855 8.005 1.48 ;
        RECT 7.145 1.095 7.285 1.48 ;
        RECT 6.316 1.225 6.456 1.48 ;
        RECT 5.305 1.225 5.445 1.48 ;
        RECT 2.835 1.24 2.975 1.48 ;
        RECT 1.505 1.24 1.645 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 8.4 0.08 ;
        RECT 7.56 -0.08 7.65 0.365 ;
        RECT 6.855 -0.08 6.995 0.26 ;
        RECT 5.95 -0.08 6.09 0.16 ;
        RECT 2.865 -0.08 3.005 0.16 ;
        RECT 1.395 -0.08 1.535 0.175 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.535 0.625 1.75 0.805 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.43 0.645 0.625 0.781 ;
        RECT 0.444 0.645 0.58 0.825 ;
        RECT 0.43 0.645 0.58 0.782 ;
        RECT 0.405 0.645 0.625 0.75 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 8.165 0.25 8.255 1.145 ;
        RECT 7.785 0.25 8.255 0.35 ;
      LAYER MET2 ;
        RECT 7.85 0.18 7.95 0.56 ;
      LAYER VIA1 ;
        RECT 7.855 0.255 7.945 0.345 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.555 0.645 7.645 1.05 ;
        RECT 7.38 0.645 7.645 0.735 ;
        RECT 7.38 0.25 7.47 0.735 ;
        RECT 7.17 0.25 7.47 0.35 ;
      LAYER MET2 ;
        RECT 7.25 0.18 7.35 0.56 ;
      LAYER VIA1 ;
        RECT 7.255 0.255 7.345 0.345 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.985 0.45 6.175 0.69 ;
      LAYER MET2 ;
        RECT 6.05 0.23 6.15 0.76 ;
      LAYER VIA1 ;
        RECT 6.055 0.455 6.145 0.545 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.715 0.74 0.805 0.906 ;
        RECT 0.646 0.896 0.761 0.951 ;
        RECT 0.684 0.861 0.715 0.99 ;
        RECT 0.281 0.915 0.684 1.005 ;
        RECT 0.225 0.825 0.35 0.972 ;
        RECT 0.225 0.715 0.315 0.972 ;
        RECT 0.271 0.915 0.684 1 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.435 1.265 0.565 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END SI
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.28 0.53 6.62 0.75 ;
      LAYER MET2 ;
        RECT 6.45 0.425 6.55 0.96 ;
      LAYER VIA1 ;
        RECT 6.455 0.655 6.545 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 7.375 1.14 7.825 1.23 ;
      RECT 7.735 0.62 7.825 1.23 ;
      RECT 6.589 1.14 7.01 1.23 ;
      RECT 6.92 0.915 7.01 1.23 ;
      RECT 5.58 1.14 6.183 1.23 ;
      RECT 6.578 1.096 6.589 1.225 ;
      RECT 5.569 1.096 5.58 1.225 ;
      RECT 4.88 1.07 4.97 1.225 ;
      RECT 6.532 1.068 6.578 1.196 ;
      RECT 5.523 1.068 5.569 1.196 ;
      RECT 4.88 1.07 5.239 1.16 ;
      RECT 4.88 1.07 5.264 1.148 ;
      RECT 7.375 0.915 7.465 1.23 ;
      RECT 6.494 1.121 6.627 1.154 ;
      RECT 6.145 1.121 6.278 1.154 ;
      RECT 6.229 1.05 6.24 1.179 ;
      RECT 5.485 1.121 5.618 1.154 ;
      RECT 6.24 1.045 6.532 1.135 ;
      RECT 5.226 1.045 5.523 1.135 ;
      RECT 6.183 1.079 6.229 1.207 ;
      RECT 5.201 1.057 5.239 1.16 ;
      RECT 6.92 0.915 7.465 1.005 ;
      RECT 7.2 0.44 7.29 1.005 ;
      RECT 7.735 0.62 8.075 0.71 ;
      RECT 6.75 0.44 7.29 0.53 ;
      RECT 6.605 0.35 6.84 0.44 ;
      RECT 6.605 0.205 6.695 0.44 ;
      RECT 6.665 0.865 6.83 1.05 ;
      RECT 6.74 0.62 6.83 1.05 ;
      RECT 5.656 0.96 6.107 1.05 ;
      RECT 4.52 0.71 4.61 1.05 ;
      RECT 5.645 0.916 5.656 1.045 ;
      RECT 5.645 0.96 6.153 1.027 ;
      RECT 5.599 0.888 5.645 1.016 ;
      RECT 6.069 0.941 6.202 0.974 ;
      RECT 6.153 0.87 6.164 0.999 ;
      RECT 5.561 0.941 5.694 0.974 ;
      RECT 6.164 0.865 6.83 0.955 ;
      RECT 5.2 0.865 5.599 0.955 ;
      RECT 6.107 0.899 6.83 0.955 ;
      RECT 5.2 0.71 5.29 0.955 ;
      RECT 4.52 0.71 5.29 0.8 ;
      RECT 6.74 0.62 7.11 0.71 ;
      RECT 4.915 0.35 5.005 0.8 ;
      RECT 4.38 0.35 5.495 0.44 ;
      RECT 3.595 0.17 3.685 0.381 ;
      RECT 5.873 0.25 6.49 0.34 ;
      RECT 5.831 0.191 5.873 0.319 ;
      RECT 5.793 0.25 6.49 0.279 ;
      RECT 3.595 0.17 5.831 0.26 ;
      RECT 3.595 0.231 5.911 0.26 ;
      RECT 5.805 0.78 6.03 0.87 ;
      RECT 5.805 0.53 5.895 0.87 ;
      RECT 5.155 0.53 5.895 0.62 ;
      RECT 5.64 0.35 5.73 0.62 ;
      RECT 5.615 0.35 5.755 0.44 ;
      RECT 3.48 1.14 4.79 1.23 ;
      RECT 4.7 0.89 4.79 1.23 ;
      RECT 3.48 1.07 3.57 1.23 ;
      RECT 4.7 0.89 5.11 0.98 ;
      RECT 3.678 0.96 4.43 1.05 ;
      RECT 4.34 0.53 4.43 1.05 ;
      RECT 3.636 0.901 3.678 1.029 ;
      RECT 3.598 0.96 4.43 0.989 ;
      RECT 2.5 0.88 3.636 0.97 ;
      RECT 2.5 0.941 3.716 0.97 ;
      RECT 2.5 0.43 2.59 0.97 ;
      RECT 4.34 0.53 4.825 0.62 ;
      RECT 2.5 0.43 3.295 0.52 ;
      RECT 3.205 0.35 3.295 0.52 ;
      RECT 3.754 0.78 4.25 0.87 ;
      RECT 4.16 0.35 4.25 0.87 ;
      RECT 3.712 0.721 3.754 0.849 ;
      RECT 3.674 0.78 4.25 0.809 ;
      RECT 2.705 0.7 3.712 0.79 ;
      RECT 2.705 0.761 3.792 0.79 ;
      RECT 3.985 0.35 4.25 0.44 ;
      RECT 1.785 0.905 1.95 0.995 ;
      RECT 1.86 0.535 1.95 0.995 ;
      RECT 3.821 0.58 4.07 0.67 ;
      RECT 3.799 0.531 3.821 0.659 ;
      RECT 3.761 0.58 4.07 0.629 ;
      RECT 3.39 0.52 3.799 0.61 ;
      RECT 3.39 0.561 3.859 0.61 ;
      RECT 1.821 0.446 1.86 0.575 ;
      RECT 1.821 0.523 1.929 0.575 ;
      RECT 1.775 0.404 1.821 0.532 ;
      RECT 1.775 0.489 1.906 0.532 ;
      RECT 3.39 0.17 3.48 0.61 ;
      RECT 1.731 0.17 1.775 0.487 ;
      RECT 1.685 0.17 1.775 0.442 ;
      RECT 2.685 0.25 3.081 0.34 ;
      RECT 2.685 0.25 3.161 0.279 ;
      RECT 3.123 0.17 3.48 0.26 ;
      RECT 3.043 0.231 3.48 0.26 ;
      RECT 3.081 0.191 3.123 0.319 ;
      RECT 1.685 0.17 2.775 0.26 ;
      RECT 3.27 1.06 3.36 1.225 ;
      RECT 2.29 1.06 3.36 1.15 ;
      RECT 2.29 0.35 2.38 1.15 ;
      RECT 2.225 0.35 2.38 0.44 ;
      RECT 1.763 1.14 2.13 1.23 ;
      RECT 2.04 0.35 2.13 1.23 ;
      RECT 1.721 1.081 1.763 1.209 ;
      RECT 1.683 1.14 2.13 1.169 ;
      RECT 0.76 1.06 1.721 1.15 ;
      RECT 0.76 1.121 1.801 1.15 ;
      RECT 1.355 0.335 1.445 1.15 ;
      RECT 1.975 0.35 2.13 0.44 ;
      RECT 1.349 0.264 1.355 0.392 ;
      RECT 1.303 0.238 1.349 0.366 ;
      RECT 1.303 0.29 1.401 0.366 ;
      RECT 1.265 0.29 1.401 0.324 ;
      RECT 0.755 0.215 1.303 0.305 ;
      RECT 0.045 1.08 0.185 1.17 ;
      RECT 0.045 0.395 0.135 1.17 ;
      RECT 1.028 0.735 1.235 0.825 ;
      RECT 1.026 0.696 1.028 0.824 ;
      RECT 0.98 0.672 1.026 0.8 ;
      RECT 0.934 0.626 0.98 0.754 ;
      RECT 0.934 0.716 1.066 0.754 ;
      RECT 0.888 0.58 0.934 0.708 ;
      RECT 0.842 0.534 0.888 0.662 ;
      RECT 0.796 0.488 0.842 0.616 ;
      RECT 0.758 0.534 0.888 0.574 ;
      RECT 0.445 0.465 0.796 0.555 ;
      RECT 0.045 0.395 0.535 0.485 ;
      RECT 0.07 0.224 0.16 0.485 ;
  END
END SDFFNSRX1H7R

MACRO SDFFNSX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNSX0P5H7R 0 0 ;
  SIZE 6.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.8 1.48 ;
        RECT 6.13 1.225 6.27 1.48 ;
        RECT 5.62 1.225 5.76 1.48 ;
        RECT 4.885 1.07 4.975 1.48 ;
        RECT 3.285 1.225 3.425 1.48 ;
        RECT 2.775 1.225 2.915 1.48 ;
        RECT 1.43 1.225 1.57 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.8 0.08 ;
        RECT 6.19 -0.08 6.28 0.345 ;
        RECT 5.685 -0.08 5.825 0.39 ;
        RECT 5.235 -0.08 5.375 0.174 ;
        RECT 2.915 -0.08 3.055 0.175 ;
        RECT 1.35 -0.08 1.49 0.175 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.55 0.625 1.75 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.62 0.595 0.815 ;
        RECT 0.425 0.62 0.595 0.75 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.425 0.262 6.575 1.15 ;
        RECT 6.395 0.262 6.575 0.352 ;
      LAYER MET2 ;
        RECT 6.45 0.425 6.55 0.96 ;
      LAYER VIA1 ;
        RECT 6.455 0.655 6.545 0.745 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.96 0.45 6.175 0.55 ;
        RECT 5.96 0.335 6.07 0.945 ;
      LAYER MET2 ;
        RECT 6.05 0.23 6.15 0.76 ;
      LAYER VIA1 ;
        RECT 6.055 0.455 6.145 0.545 ;
    END
  END QN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.905 0.82 0.995 ;
        RECT 0.73 0.74 0.82 0.995 ;
        RECT 0.225 0.825 0.35 0.995 ;
        RECT 0.225 0.615 0.315 0.995 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.185 0.455 1.275 0.605 ;
        RECT 1.05 0.455 1.275 0.575 ;
        RECT 1.025 0.425 1.15 0.545 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END SI
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.005 0.65 5.195 0.795 ;
      LAYER MET2 ;
        RECT 5.05 0.43 5.15 0.96 ;
      LAYER VIA1 ;
        RECT 5.055 0.655 5.145 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 5.355 1.035 6.329 1.125 ;
      RECT 6.239 0.62 6.329 1.125 ;
      RECT 5.72 0.48 5.81 1.125 ;
      RECT 4.865 0.435 4.955 0.575 ;
      RECT 5.293 0.48 5.81 0.57 ;
      RECT 4.865 0.47 5.575 0.56 ;
      RECT 5.435 0.375 5.575 0.57 ;
      RECT 5.15 0.89 5.24 1.195 ;
      RECT 3.98 1.085 4.775 1.175 ;
      RECT 4.685 0.35 4.775 1.175 ;
      RECT 4.685 0.89 5.274 0.98 ;
      RECT 4.685 0.89 5.331 0.946 ;
      RECT 5.285 0.66 5.375 0.901 ;
      RECT 5.236 0.888 5.375 0.901 ;
      RECT 5.274 0.846 5.285 0.975 ;
      RECT 5.24 0.869 5.375 0.901 ;
      RECT 5.285 0.66 5.63 0.75 ;
      RECT 4.48 0.35 4.775 0.44 ;
      RECT 4.995 0.17 5.085 0.35 ;
      RECT 3.65 0.17 5.085 0.26 ;
      RECT 2.745 1.045 3.8 1.135 ;
      RECT 3.71 0.905 3.8 1.135 ;
      RECT 2.745 0.86 2.835 1.135 ;
      RECT 3.71 0.905 4.595 0.995 ;
      RECT 4.505 0.53 4.595 0.995 ;
      RECT 4.285 0.53 4.595 0.62 ;
      RECT 4.285 0.35 4.375 0.62 ;
      RECT 4.2 0.35 4.375 0.44 ;
      RECT 3.105 0.865 3.61 0.955 ;
      RECT 3.52 0.582 3.61 0.955 ;
      RECT 3.52 0.725 4.415 0.815 ;
      RECT 2.385 0.563 2.475 0.745 ;
      RECT 3.755 0.69 3.895 0.815 ;
      RECT 3.481 0.494 3.52 0.623 ;
      RECT 2.385 0.563 2.534 0.584 ;
      RECT 3.443 0.537 3.566 0.584 ;
      RECT 2.496 0.475 3.481 0.565 ;
      RECT 2.475 0.485 2.496 0.614 ;
      RECT 2.431 0.518 3.52 0.565 ;
      RECT 3.245 0.385 3.385 0.565 ;
      RECT 1.74 0.915 1.935 1.005 ;
      RECT 1.845 0.17 1.935 1.005 ;
      RECT 3.99 0.525 4.165 0.615 ;
      RECT 3.99 0.365 4.08 0.615 ;
      RECT 3.589 0.365 4.08 0.455 ;
      RECT 3.56 0.312 3.589 0.441 ;
      RECT 1.68 0.28 1.935 0.37 ;
      RECT 3.516 0.346 3.627 0.404 ;
      RECT 3.47 0.185 3.56 0.359 ;
      RECT 2.716 0.265 3.131 0.355 ;
      RECT 2.705 0.221 2.716 0.35 ;
      RECT 2.659 0.193 2.705 0.321 ;
      RECT 2.659 0.265 3.211 0.294 ;
      RECT 3.173 0.185 3.56 0.275 ;
      RECT 3.093 0.246 3.56 0.275 ;
      RECT 3.131 0.206 3.173 0.334 ;
      RECT 2.621 0.246 2.754 0.279 ;
      RECT 1.845 0.17 2.659 0.26 ;
      RECT 2.275 0.9 2.365 1.195 ;
      RECT 2.205 0.9 2.489 0.99 ;
      RECT 2.205 0.9 2.535 0.967 ;
      RECT 2.451 0.881 2.565 0.929 ;
      RECT 2.205 0.36 2.295 0.99 ;
      RECT 2.489 0.839 2.611 0.891 ;
      RECT 2.535 0.801 2.565 0.929 ;
      RECT 2.565 0.68 2.655 0.846 ;
      RECT 3.285 0.68 3.425 0.775 ;
      RECT 2.565 0.68 3.425 0.77 ;
      RECT 2.205 0.36 2.39 0.45 ;
      RECT 1.706 1.14 2.115 1.23 ;
      RECT 2.025 0.35 2.115 1.23 ;
      RECT 1.695 1.096 1.706 1.225 ;
      RECT 1.649 1.068 1.695 1.196 ;
      RECT 1.611 1.121 1.744 1.154 ;
      RECT 0.925 1.045 1.649 1.135 ;
      RECT 1.37 0.275 1.46 1.135 ;
      RECT 1.247 0.275 1.46 0.365 ;
      RECT 1.225 0.226 1.247 0.354 ;
      RECT 1.187 0.275 1.46 0.324 ;
      RECT 0.755 0.215 1.225 0.305 ;
      RECT 0.755 0.256 1.285 0.305 ;
      RECT 0.045 1.08 0.185 1.17 ;
      RECT 0.045 0.255 0.135 1.17 ;
      RECT 0.93 0.74 1.225 0.83 ;
      RECT 0.93 0.68 1.02 0.83 ;
      RECT 0.908 0.572 0.93 0.7 ;
      RECT 0.908 0.65 1.019 0.7 ;
      RECT 0.862 0.538 0.908 0.666 ;
      RECT 0.862 0.606 0.976 0.666 ;
      RECT 0.824 0.515 0.862 0.624 ;
      RECT 0.7 0.515 0.862 0.605 ;
      RECT 0.7 0.395 0.79 0.605 ;
      RECT 0.045 0.395 0.79 0.485 ;
      RECT 0.045 0.255 0.16 0.485 ;
  END
END SDFFNSX0P5H7R

MACRO SDFFNSX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNSX1H7R 0 0 ;
  SIZE 6.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.8 1.48 ;
        RECT 6.13 1.225 6.27 1.48 ;
        RECT 5.62 1.225 5.76 1.48 ;
        RECT 4.885 1.07 4.975 1.48 ;
        RECT 3.285 1.225 3.425 1.48 ;
        RECT 2.775 1.225 2.915 1.48 ;
        RECT 1.43 1.225 1.57 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.8 0.08 ;
        RECT 6.19 -0.08 6.28 0.345 ;
        RECT 5.685 -0.08 5.825 0.38 ;
        RECT 5.235 -0.08 5.375 0.174 ;
        RECT 2.915 -0.08 3.055 0.175 ;
        RECT 1.35 -0.08 1.49 0.175 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.55 0.625 1.75 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.62 0.595 0.815 ;
        RECT 0.425 0.62 0.595 0.75 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.425 0.305 6.575 1.15 ;
        RECT 6.385 0.305 6.575 0.395 ;
      LAYER MET2 ;
        RECT 6.45 0.425 6.55 0.96 ;
      LAYER VIA1 ;
        RECT 6.455 0.655 6.545 0.745 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.96 0.45 6.175 0.55 ;
        RECT 5.96 0.335 6.07 0.945 ;
      LAYER MET2 ;
        RECT 6.05 0.23 6.15 0.76 ;
      LAYER VIA1 ;
        RECT 6.055 0.455 6.145 0.545 ;
    END
  END QN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.905 0.82 0.995 ;
        RECT 0.73 0.74 0.82 0.995 ;
        RECT 0.225 0.825 0.35 0.995 ;
        RECT 0.225 0.615 0.315 0.995 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.185 0.455 1.275 0.605 ;
        RECT 1.05 0.455 1.275 0.575 ;
        RECT 1.02 0.425 1.15 0.545 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END SI
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.005 0.65 5.195 0.795 ;
      LAYER MET2 ;
        RECT 5.05 0.43 5.15 0.96 ;
      LAYER VIA1 ;
        RECT 5.055 0.655 5.145 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 5.355 1.035 6.329 1.125 ;
      RECT 6.239 0.62 6.329 1.125 ;
      RECT 5.72 0.47 5.81 1.125 ;
      RECT 4.865 0.435 4.955 0.575 ;
      RECT 4.865 0.47 5.81 0.56 ;
      RECT 5.435 0.375 5.575 0.56 ;
      RECT 5.15 0.89 5.24 1.195 ;
      RECT 3.98 1.085 4.775 1.175 ;
      RECT 4.685 0.35 4.775 1.175 ;
      RECT 4.685 0.89 5.274 0.98 ;
      RECT 4.685 0.89 5.331 0.946 ;
      RECT 5.285 0.66 5.375 0.901 ;
      RECT 5.236 0.888 5.375 0.901 ;
      RECT 5.274 0.846 5.285 0.975 ;
      RECT 5.24 0.869 5.375 0.901 ;
      RECT 5.285 0.66 5.63 0.75 ;
      RECT 4.48 0.35 4.775 0.44 ;
      RECT 4.995 0.17 5.085 0.35 ;
      RECT 3.65 0.17 5.085 0.26 ;
      RECT 2.745 1.045 3.8 1.135 ;
      RECT 3.71 0.905 3.8 1.135 ;
      RECT 2.745 0.86 2.835 1.135 ;
      RECT 3.71 0.905 4.595 0.995 ;
      RECT 4.505 0.53 4.595 0.995 ;
      RECT 4.285 0.53 4.595 0.62 ;
      RECT 4.285 0.35 4.375 0.62 ;
      RECT 4.2 0.35 4.375 0.44 ;
      RECT 3.105 0.865 3.61 0.955 ;
      RECT 3.52 0.582 3.61 0.955 ;
      RECT 3.52 0.725 4.415 0.815 ;
      RECT 2.385 0.563 2.475 0.745 ;
      RECT 3.52 0.705 4.255 0.815 ;
      RECT 3.481 0.494 3.52 0.623 ;
      RECT 2.385 0.563 2.534 0.584 ;
      RECT 3.443 0.537 3.566 0.584 ;
      RECT 2.496 0.475 3.481 0.565 ;
      RECT 2.475 0.485 2.496 0.614 ;
      RECT 2.431 0.518 3.52 0.565 ;
      RECT 3.245 0.385 3.385 0.565 ;
      RECT 1.74 0.915 1.935 1.005 ;
      RECT 1.845 0.17 1.935 1.005 ;
      RECT 3.99 0.525 4.165 0.615 ;
      RECT 3.99 0.365 4.08 0.615 ;
      RECT 3.589 0.365 4.08 0.455 ;
      RECT 3.56 0.312 3.589 0.441 ;
      RECT 1.68 0.28 1.935 0.37 ;
      RECT 3.516 0.346 3.627 0.404 ;
      RECT 3.47 0.185 3.56 0.359 ;
      RECT 2.716 0.265 3.131 0.355 ;
      RECT 2.705 0.221 2.716 0.35 ;
      RECT 2.659 0.193 2.705 0.321 ;
      RECT 2.659 0.265 3.211 0.294 ;
      RECT 3.173 0.185 3.56 0.275 ;
      RECT 3.093 0.246 3.56 0.275 ;
      RECT 3.131 0.206 3.173 0.334 ;
      RECT 2.621 0.246 2.754 0.279 ;
      RECT 1.845 0.17 2.659 0.26 ;
      RECT 2.205 0.9 2.365 1.195 ;
      RECT 2.205 0.9 2.489 0.99 ;
      RECT 2.205 0.9 2.535 0.967 ;
      RECT 2.451 0.881 2.565 0.929 ;
      RECT 2.205 0.36 2.295 1.195 ;
      RECT 2.489 0.839 2.611 0.891 ;
      RECT 2.535 0.801 2.565 0.929 ;
      RECT 2.565 0.68 2.655 0.846 ;
      RECT 3.285 0.68 3.425 0.775 ;
      RECT 2.565 0.68 3.425 0.77 ;
      RECT 2.205 0.36 2.39 0.45 ;
      RECT 1.706 1.14 2.115 1.23 ;
      RECT 2.025 0.35 2.115 1.23 ;
      RECT 1.695 1.096 1.706 1.225 ;
      RECT 1.649 1.068 1.695 1.196 ;
      RECT 1.611 1.121 1.744 1.154 ;
      RECT 0.925 1.045 1.649 1.135 ;
      RECT 1.37 0.275 1.46 1.135 ;
      RECT 1.247 0.275 1.46 0.365 ;
      RECT 1.225 0.226 1.247 0.354 ;
      RECT 1.187 0.275 1.46 0.324 ;
      RECT 0.755 0.215 1.225 0.305 ;
      RECT 0.755 0.256 1.285 0.305 ;
      RECT 0.045 1.08 0.185 1.17 ;
      RECT 0.045 0.255 0.135 1.17 ;
      RECT 0.93 0.74 1.225 0.83 ;
      RECT 0.93 0.68 1.02 0.83 ;
      RECT 0.908 0.572 0.93 0.7 ;
      RECT 0.908 0.65 1.019 0.7 ;
      RECT 0.862 0.538 0.908 0.666 ;
      RECT 0.862 0.606 0.976 0.666 ;
      RECT 0.824 0.515 0.862 0.624 ;
      RECT 0.7 0.515 0.862 0.605 ;
      RECT 0.7 0.395 0.79 0.605 ;
      RECT 0.045 0.395 0.79 0.485 ;
      RECT 0.045 0.255 0.16 0.485 ;
  END
END SDFFNSX1H7R

MACRO SDFFNSX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNSX2H7R 0 0 ;
  SIZE 6.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.8 1.48 ;
        RECT 6.13 1.225 6.27 1.48 ;
        RECT 5.62 1.225 5.76 1.48 ;
        RECT 4.885 1.07 4.975 1.48 ;
        RECT 3.285 1.225 3.425 1.48 ;
        RECT 2.775 1.225 2.915 1.48 ;
        RECT 1.43 1.225 1.57 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.8 0.08 ;
        RECT 6.19 -0.08 6.28 0.345 ;
        RECT 5.685 -0.08 5.825 0.35 ;
        RECT 5.235 -0.08 5.375 0.174 ;
        RECT 2.915 -0.08 3.055 0.175 ;
        RECT 1.35 -0.08 1.49 0.175 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.55 0.625 1.75 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.62 0.595 0.815 ;
        RECT 0.425 0.62 0.595 0.75 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.425 0.305 6.575 1.15 ;
        RECT 6.39 0.305 6.575 0.395 ;
      LAYER MET2 ;
        RECT 6.45 0.425 6.55 0.96 ;
      LAYER VIA1 ;
        RECT 6.455 0.655 6.545 0.745 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.96 0.45 6.175 0.55 ;
        RECT 5.96 0.335 6.07 0.945 ;
      LAYER MET2 ;
        RECT 6.05 0.23 6.15 0.76 ;
      LAYER VIA1 ;
        RECT 6.055 0.455 6.145 0.545 ;
    END
  END QN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.905 0.82 0.995 ;
        RECT 0.73 0.74 0.82 0.995 ;
        RECT 0.225 0.825 0.35 0.995 ;
        RECT 0.225 0.615 0.315 0.995 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.185 0.455 1.275 0.605 ;
        RECT 1.05 0.455 1.275 0.575 ;
        RECT 1.02 0.425 1.15 0.545 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END SI
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.005 0.65 5.195 0.795 ;
      LAYER MET2 ;
        RECT 5.05 0.43 5.15 0.96 ;
      LAYER VIA1 ;
        RECT 5.055 0.655 5.145 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 5.355 1.035 6.329 1.125 ;
      RECT 6.239 0.62 6.329 1.125 ;
      RECT 5.72 0.47 5.81 1.125 ;
      RECT 4.865 0.435 4.955 0.575 ;
      RECT 4.865 0.47 5.81 0.56 ;
      RECT 5.435 0.375 5.575 0.56 ;
      RECT 5.15 0.89 5.24 1.195 ;
      RECT 3.98 1.085 4.775 1.175 ;
      RECT 4.685 0.35 4.775 1.175 ;
      RECT 4.685 0.89 5.274 0.98 ;
      RECT 4.685 0.89 5.331 0.946 ;
      RECT 5.285 0.66 5.375 0.901 ;
      RECT 5.236 0.888 5.375 0.901 ;
      RECT 5.274 0.846 5.285 0.975 ;
      RECT 5.24 0.869 5.375 0.901 ;
      RECT 5.285 0.66 5.63 0.75 ;
      RECT 4.48 0.35 4.775 0.44 ;
      RECT 4.995 0.17 5.085 0.35 ;
      RECT 3.65 0.17 5.085 0.26 ;
      RECT 2.745 1.045 3.8 1.135 ;
      RECT 3.71 0.905 3.8 1.135 ;
      RECT 2.745 0.86 2.835 1.135 ;
      RECT 3.71 0.905 4.595 0.995 ;
      RECT 4.505 0.53 4.595 0.995 ;
      RECT 4.285 0.53 4.595 0.62 ;
      RECT 4.285 0.35 4.375 0.62 ;
      RECT 4.2 0.35 4.375 0.44 ;
      RECT 3.105 0.865 3.61 0.955 ;
      RECT 3.52 0.582 3.61 0.955 ;
      RECT 3.52 0.725 4.415 0.815 ;
      RECT 2.385 0.563 2.475 0.745 ;
      RECT 3.52 0.705 3.895 0.815 ;
      RECT 3.481 0.494 3.52 0.623 ;
      RECT 2.385 0.563 2.534 0.584 ;
      RECT 3.443 0.537 3.566 0.584 ;
      RECT 2.496 0.475 3.481 0.565 ;
      RECT 2.475 0.485 2.496 0.614 ;
      RECT 2.431 0.518 3.52 0.565 ;
      RECT 3.245 0.385 3.385 0.565 ;
      RECT 1.74 0.915 1.935 1.005 ;
      RECT 1.845 0.17 1.935 1.005 ;
      RECT 3.99 0.525 4.165 0.615 ;
      RECT 3.99 0.365 4.08 0.615 ;
      RECT 3.589 0.365 4.08 0.455 ;
      RECT 3.56 0.312 3.589 0.441 ;
      RECT 1.68 0.28 1.935 0.37 ;
      RECT 3.516 0.346 3.627 0.404 ;
      RECT 3.47 0.185 3.56 0.359 ;
      RECT 2.716 0.265 3.131 0.355 ;
      RECT 2.705 0.221 2.716 0.35 ;
      RECT 2.659 0.193 2.705 0.321 ;
      RECT 2.659 0.265 3.211 0.294 ;
      RECT 3.173 0.185 3.56 0.275 ;
      RECT 3.093 0.246 3.56 0.275 ;
      RECT 3.131 0.206 3.173 0.334 ;
      RECT 2.621 0.246 2.754 0.279 ;
      RECT 1.845 0.17 2.659 0.26 ;
      RECT 2.275 0.9 2.365 1.195 ;
      RECT 2.205 0.9 2.489 0.99 ;
      RECT 2.205 0.9 2.535 0.967 ;
      RECT 2.451 0.881 2.565 0.929 ;
      RECT 2.205 0.36 2.295 0.99 ;
      RECT 2.489 0.839 2.611 0.891 ;
      RECT 2.535 0.801 2.565 0.929 ;
      RECT 2.565 0.68 2.655 0.846 ;
      RECT 3.285 0.68 3.425 0.775 ;
      RECT 2.565 0.68 3.425 0.77 ;
      RECT 2.205 0.36 2.39 0.45 ;
      RECT 1.706 1.14 2.115 1.23 ;
      RECT 2.025 0.35 2.115 1.23 ;
      RECT 1.695 1.096 1.706 1.225 ;
      RECT 1.649 1.068 1.695 1.196 ;
      RECT 1.611 1.121 1.744 1.154 ;
      RECT 0.925 1.045 1.649 1.135 ;
      RECT 1.37 0.275 1.46 1.135 ;
      RECT 1.247 0.275 1.46 0.365 ;
      RECT 1.225 0.226 1.247 0.354 ;
      RECT 1.187 0.275 1.46 0.324 ;
      RECT 0.755 0.215 1.225 0.305 ;
      RECT 0.755 0.256 1.285 0.305 ;
      RECT 0.045 1.08 0.185 1.17 ;
      RECT 0.045 0.255 0.135 1.17 ;
      RECT 0.93 0.74 1.225 0.83 ;
      RECT 0.93 0.68 1.02 0.83 ;
      RECT 0.908 0.572 0.93 0.7 ;
      RECT 0.908 0.65 1.019 0.7 ;
      RECT 0.862 0.538 0.908 0.666 ;
      RECT 0.862 0.606 0.976 0.666 ;
      RECT 0.824 0.515 0.862 0.624 ;
      RECT 0.7 0.515 0.862 0.605 ;
      RECT 0.7 0.395 0.79 0.605 ;
      RECT 0.045 0.395 0.79 0.485 ;
      RECT 0.045 0.255 0.16 0.485 ;
  END
END SDFFNSX2H7R

MACRO SDFFNX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNX0P5H7R 0 0 ;
  SIZE 6.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.8 1.48 ;
        RECT 6.31 1.035 6.4 1.48 ;
        RECT 5.59 1.05 5.68 1.48 ;
        RECT 4.795 1.08 4.935 1.48 ;
        RECT 3.525 1.24 3.665 1.48 ;
        RECT 2.6 1.24 2.74 1.48 ;
        RECT 1.145 1.24 1.285 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.8 0.08 ;
        RECT 6.31 -0.08 6.4 0.345 ;
        RECT 5.805 -0.08 5.895 0.33 ;
        RECT 4.795 -0.08 4.935 0.19 ;
        RECT 3.535 -0.08 3.675 0.16 ;
        RECT 2.59 -0.08 2.73 0.16 ;
        RECT 1.08 -0.08 1.22 0.16 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.22 0.65 3.49 0.75 ;
      LAYER MET2 ;
        RECT 3.25 0.43 3.35 0.96 ;
      LAYER VIA1 ;
        RECT 3.255 0.655 3.345 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.95 0.466 6.16 0.556 ;
        RECT 6.055 0.225 6.16 0.556 ;
        RECT 5.95 0.466 6.04 1.045 ;
      LAYER MET2 ;
        RECT 6.05 0.18 6.15 0.56 ;
      LAYER VIA1 ;
        RECT 6.055 0.255 6.145 0.345 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.585 0.255 6.745 1.045 ;
      LAYER MET2 ;
        RECT 6.65 0.425 6.75 0.96 ;
      LAYER VIA1 ;
        RECT 6.655 0.655 6.745 0.745 ;
    END
  END QN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.285 0.508 1.375 0.665 ;
        RECT 0.66 0.478 1.36 0.545 ;
        RECT 0.66 0.455 1.314 0.545 ;
        RECT 1.276 0.508 1.375 0.55 ;
        RECT 0.66 0.455 0.75 0.605 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1 0.64 1.18 0.79 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.77 1.135 6.22 1.225 ;
      RECT 6.13 0.685 6.22 1.225 ;
      RECT 5.77 0.71 5.86 1.225 ;
      RECT 5.34 0.71 5.43 1.045 ;
      RECT 4.615 0.71 5.86 0.8 ;
      RECT 6.13 0.685 6.49 0.775 ;
      RECT 5.54 0.31 5.63 0.8 ;
      RECT 4.2 0.28 4.29 1.03 ;
      RECT 4.2 0.28 5.014 0.37 ;
      RECT 4.2 0.28 5.06 0.347 ;
      RECT 4.976 0.261 5.086 0.311 ;
      RECT 5.014 0.219 5.124 0.279 ;
      RECT 5.06 0.183 5.086 0.311 ;
      RECT 5.086 0.17 5.46 0.26 ;
      RECT 2.83 1.14 3.32 1.23 ;
      RECT 1.875 1.14 2.4 1.23 ;
      RECT 4.02 1.12 4.47 1.21 ;
      RECT 4.38 0.46 4.47 1.21 ;
      RECT 3.23 1.06 4.11 1.15 ;
      RECT 2.31 1.06 2.92 1.15 ;
      RECT 1.875 0.505 1.965 1.23 ;
      RECT 4.02 0.72 4.11 1.21 ;
      RECT 4.38 0.9 5.225 0.99 ;
      RECT 4.38 0.46 5.255 0.55 ;
      RECT 5.165 0.35 5.255 0.55 ;
      RECT 5.165 0.35 5.305 0.44 ;
      RECT 3.23 0.88 3.93 0.97 ;
      RECT 3.84 0.29 3.93 0.97 ;
      RECT 3.84 0.475 4.04 0.615 ;
      RECT 2.235 0.25 2.325 0.575 ;
      RECT 3.27 0.29 3.93 0.38 ;
      RECT 2.235 0.25 2.91 0.34 ;
      RECT 3.27 0.17 3.36 0.38 ;
      RECT 2.82 0.17 3.36 0.26 ;
      RECT 3.025 0.35 3.115 1.05 ;
      RECT 3.66 0.47 3.75 0.61 ;
      RECT 2.44 0.51 3.115 0.6 ;
      RECT 3 0.47 3.75 0.56 ;
      RECT 3 0.35 3.14 0.56 ;
      RECT 2.055 0.27 2.145 1.05 ;
      RECT 2.055 0.74 2.92 0.83 ;
      RECT 0.635 1.06 1.785 1.15 ;
      RECT 1.695 0.17 1.785 1.15 ;
      RECT 1.695 0.17 1.825 0.37 ;
      RECT 0.535 0.25 1.299 0.34 ;
      RECT 0.535 0.25 1.379 0.279 ;
      RECT 1.341 0.17 1.825 0.26 ;
      RECT 1.261 0.231 1.825 0.26 ;
      RECT 1.299 0.191 1.341 0.319 ;
      RECT 0.81 0.88 1.58 0.97 ;
      RECT 1.49 0.35 1.58 0.97 ;
      RECT 0.81 0.695 0.9 0.97 ;
      RECT 0.4 0.695 0.9 0.785 ;
      RECT 0.4 0.465 0.49 0.785 ;
      RECT 1.44 0.35 1.58 0.44 ;
  END
END SDFFNX0P5H7R

MACRO SDFFNX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNX1H7R 0 0 ;
  SIZE 6.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.8 1.48 ;
        RECT 6.335 1.03 6.425 1.48 ;
        RECT 5.59 1.05 5.68 1.48 ;
        RECT 4.795 1.11 4.935 1.48 ;
        RECT 3.525 1.24 3.665 1.48 ;
        RECT 2.6 1.095 2.74 1.48 ;
        RECT 1.145 1.24 1.285 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.8 0.08 ;
        RECT 6.335 -0.08 6.425 0.345 ;
        RECT 5.825 -0.08 5.915 0.36 ;
        RECT 4.795 -0.08 4.935 0.16 ;
        RECT 3.535 -0.08 3.675 0.2 ;
        RECT 2.59 -0.08 2.73 0.27 ;
        RECT 1.095 -0.08 1.235 0.16 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.22 0.65 3.445 0.77 ;
      LAYER MET2 ;
        RECT 3.25 0.43 3.35 0.96 ;
      LAYER VIA1 ;
        RECT 3.255 0.655 3.345 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.95 0.455 6.175 0.545 ;
        RECT 6.085 0.295 6.175 0.545 ;
        RECT 5.95 0.455 6.04 0.985 ;
      LAYER MET2 ;
        RECT 6.05 0.23 6.15 0.76 ;
      LAYER VIA1 ;
        RECT 6.055 0.455 6.145 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.61 0.295 6.745 0.985 ;
      LAYER MET2 ;
        RECT 6.65 0.425 6.75 0.96 ;
      LAYER VIA1 ;
        RECT 6.655 0.655 6.745 0.745 ;
    END
  END QN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.285 0.455 1.375 0.605 ;
        RECT 0.67 0.455 1.375 0.545 ;
        RECT 0.67 0.455 0.76 0.605 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1 0.64 1.18 0.79 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.77 1.075 6.22 1.165 ;
      RECT 6.13 0.685 6.22 1.165 ;
      RECT 5.77 0.71 5.86 1.165 ;
      RECT 5.34 0.71 5.43 1.045 ;
      RECT 4.615 0.71 5.86 0.8 ;
      RECT 6.13 0.685 6.515 0.775 ;
      RECT 5.55 0.35 5.64 0.8 ;
      RECT 5.5 0.35 5.64 0.44 ;
      RECT 4.2 0.28 4.29 1.025 ;
      RECT 4.2 0.28 4.984 0.37 ;
      RECT 4.2 0.28 5.03 0.347 ;
      RECT 4.946 0.261 5.056 0.311 ;
      RECT 4.984 0.219 5.094 0.279 ;
      RECT 5.03 0.183 5.056 0.311 ;
      RECT 5.056 0.17 5.46 0.26 ;
      RECT 2.83 1.14 3.32 1.23 ;
      RECT 1.875 1.14 2.4 1.23 ;
      RECT 2.31 0.915 2.4 1.23 ;
      RECT 4.02 1.115 4.525 1.205 ;
      RECT 4.435 0.46 4.525 1.205 ;
      RECT 3.23 1.06 4.11 1.15 ;
      RECT 2.83 0.915 2.92 1.23 ;
      RECT 1.875 0.485 1.965 1.23 ;
      RECT 4.02 0.69 4.11 1.205 ;
      RECT 4.435 0.93 5.225 1.02 ;
      RECT 2.31 0.915 2.92 1.005 ;
      RECT 4.435 0.46 5.225 0.55 ;
      RECT 5.135 0.35 5.225 0.55 ;
      RECT 5.135 0.35 5.275 0.44 ;
      RECT 3.23 0.88 3.93 0.97 ;
      RECT 3.84 0.29 3.93 0.97 ;
      RECT 2.235 0.36 2.325 0.625 ;
      RECT 3.84 0.46 4.04 0.6 ;
      RECT 2.235 0.36 2.91 0.45 ;
      RECT 2.82 0.17 2.91 0.45 ;
      RECT 3.27 0.29 3.93 0.38 ;
      RECT 3.27 0.17 3.36 0.38 ;
      RECT 2.82 0.17 3.36 0.26 ;
      RECT 3.025 0.35 3.115 1.05 ;
      RECT 2.46 0.54 3.115 0.63 ;
      RECT 3.66 0.47 3.75 0.62 ;
      RECT 3 0.47 3.75 0.56 ;
      RECT 3 0.35 3.14 0.56 ;
      RECT 2.055 0.27 2.145 1.05 ;
      RECT 2.055 0.72 2.92 0.81 ;
      RECT 0.635 1.06 1.785 1.15 ;
      RECT 1.695 0.17 1.785 1.15 ;
      RECT 1.695 0.17 1.825 0.365 ;
      RECT 0.505 0.25 1.339 0.34 ;
      RECT 0.505 0.25 1.419 0.279 ;
      RECT 1.381 0.17 1.825 0.26 ;
      RECT 1.301 0.231 1.825 0.26 ;
      RECT 1.339 0.191 1.381 0.319 ;
      RECT 0.81 0.88 1.605 0.97 ;
      RECT 1.515 0.35 1.605 0.97 ;
      RECT 0.81 0.725 0.9 0.97 ;
      RECT 0.4 0.725 0.9 0.815 ;
      RECT 0.4 0.465 0.49 0.815 ;
      RECT 1.465 0.35 1.605 0.44 ;
  END
END SDFFNX1H7R

MACRO SDFFNX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNX2H7R 0 0 ;
  SIZE 7 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7 1.48 ;
        RECT 6.38 1.055 6.47 1.48 ;
        RECT 5.59 1.07 5.68 1.48 ;
        RECT 4.795 1.05 4.935 1.48 ;
        RECT 3.525 1.24 3.665 1.48 ;
        RECT 2.6 1.24 2.74 1.48 ;
        RECT 1.145 1.24 1.285 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7 0.08 ;
        RECT 6.38 -0.08 6.47 0.345 ;
        RECT 5.815 -0.08 5.905 0.35 ;
        RECT 4.795 -0.08 4.935 0.16 ;
        RECT 3.535 -0.08 3.645 0.2 ;
        RECT 2.59 -0.08 2.73 0.24 ;
        RECT 1.055 -0.08 1.195 0.185 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.225 0.65 3.495 0.75 ;
      LAYER MET2 ;
        RECT 3.25 0.43 3.35 0.96 ;
      LAYER VIA1 ;
        RECT 3.255 0.655 3.345 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.965 0.455 6.175 0.545 ;
        RECT 6.085 0.335 6.175 0.545 ;
        RECT 5.965 0.455 6.055 0.945 ;
      LAYER MET2 ;
        RECT 6.05 0.23 6.15 0.76 ;
      LAYER VIA1 ;
        RECT 6.055 0.455 6.145 0.545 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.655 0.28 6.75 0.945 ;
      LAYER MET2 ;
        RECT 6.65 0.425 6.75 0.96 ;
      LAYER VIA1 ;
        RECT 6.655 0.655 6.745 0.745 ;
    END
  END QN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.285 0.455 1.375 0.63 ;
        RECT 0.66 0.455 1.375 0.545 ;
        RECT 0.66 0.455 0.75 0.605 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1 0.64 1.18 0.79 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.77 1.035 6.29 1.125 ;
      RECT 6.2 0.645 6.29 1.125 ;
      RECT 5.34 0.675 5.43 1.065 ;
      RECT 5.77 0.675 5.86 1.125 ;
      RECT 4.645 0.675 5.86 0.765 ;
      RECT 6.2 0.645 6.565 0.735 ;
      RECT 5.555 0.275 5.645 0.765 ;
      RECT 4.225 0.25 4.315 0.97 ;
      RECT 4.225 0.25 5.014 0.34 ;
      RECT 4.225 0.25 5.094 0.279 ;
      RECT 5.056 0.17 5.46 0.26 ;
      RECT 4.976 0.231 5.46 0.26 ;
      RECT 5.014 0.191 5.056 0.319 ;
      RECT 4.02 1.14 4.495 1.23 ;
      RECT 4.405 0.46 4.495 1.23 ;
      RECT 1.875 1.14 2.4 1.23 ;
      RECT 2.83 1.095 3.32 1.185 ;
      RECT 3.23 1.06 4.11 1.15 ;
      RECT 2.31 1.06 2.92 1.15 ;
      RECT 1.875 0.505 1.965 1.23 ;
      RECT 4.405 0.87 5.225 0.96 ;
      RECT 4.405 0.46 5.225 0.55 ;
      RECT 5.135 0.35 5.225 0.55 ;
      RECT 5.135 0.35 5.275 0.44 ;
      RECT 3.23 0.88 3.93 0.97 ;
      RECT 3.84 0.17 3.93 0.97 ;
      RECT 2.255 0.33 2.345 0.6 ;
      RECT 2.255 0.33 2.91 0.42 ;
      RECT 2.82 0.17 2.91 0.42 ;
      RECT 3.27 0.29 3.93 0.38 ;
      RECT 3.27 0.17 3.36 0.38 ;
      RECT 3.84 0.17 4.08 0.26 ;
      RECT 2.82 0.17 3.36 0.26 ;
      RECT 3 0.35 3.115 1.005 ;
      RECT 3.66 0.47 3.75 0.64 ;
      RECT 2.46 0.51 3.115 0.6 ;
      RECT 3 0.47 3.75 0.56 ;
      RECT 3 0.35 3.14 0.56 ;
      RECT 2.075 0.29 2.165 1.05 ;
      RECT 2.075 0.705 2.89 0.795 ;
      RECT 0.635 1.06 1.785 1.15 ;
      RECT 1.695 0.17 1.785 1.15 ;
      RECT 1.695 0.17 1.825 0.365 ;
      RECT 0.535 0.275 1.375 0.365 ;
      RECT 1.285 0.17 1.375 0.365 ;
      RECT 1.285 0.17 1.825 0.26 ;
      RECT 0.81 0.88 1.605 0.97 ;
      RECT 1.515 0.35 1.605 0.97 ;
      RECT 0.81 0.725 0.9 0.97 ;
      RECT 0.4 0.725 0.9 0.815 ;
      RECT 0.4 0.485 0.49 0.815 ;
      RECT 1.465 0.35 1.605 0.44 ;
  END
END SDFFNX2H7R

MACRO SDFFNX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNX3H7R 0 0 ;
  SIZE 7.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7.4 1.48 ;
        RECT 6.895 1.07 6.985 1.48 ;
        RECT 6.415 1.04 6.505 1.48 ;
        RECT 5.69 1.04 5.78 1.48 ;
        RECT 4.895 1.11 5.035 1.48 ;
        RECT 3.625 1.24 3.765 1.48 ;
        RECT 2.7 1.24 2.84 1.48 ;
        RECT 1.24 1.24 1.38 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7.4 0.08 ;
        RECT 6.895 -0.08 6.985 0.33 ;
        RECT 6.405 -0.08 6.495 0.37 ;
        RECT 5.905 -0.08 5.995 0.35 ;
        RECT 4.895 -0.08 5.035 0.16 ;
        RECT 3.635 -0.08 3.745 0.2 ;
        RECT 2.69 -0.08 2.83 0.16 ;
        RECT 1.14 -0.08 1.28 0.16 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.37 0.65 3.595 0.77 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.26 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.055 0.455 6.245 0.545 ;
        RECT 6.155 0.29 6.245 0.545 ;
        RECT 6.055 0.455 6.145 1.05 ;
      LAYER MET2 ;
        RECT 6.05 0.43 6.15 0.96 ;
      LAYER VIA1 ;
        RECT 6.055 0.655 6.145 0.745 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.145 0.26 7.235 1.045 ;
        RECT 6.645 0.855 7.235 0.945 ;
        RECT 6.635 0.42 7.235 0.51 ;
        RECT 6.645 0.855 6.735 1.045 ;
        RECT 6.635 0.245 6.725 0.51 ;
      LAYER MET2 ;
        RECT 7.05 0.63 7.15 1.16 ;
      LAYER VIA1 ;
        RECT 7.055 0.855 7.145 0.945 ;
    END
  END QN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.365 0.43 1.455 0.755 ;
        RECT 0.655 0.43 1.455 0.52 ;
        RECT 0.655 0.425 0.81 0.605 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.625 1.235 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.875 1.14 6.325 1.23 ;
      RECT 6.235 0.675 6.325 1.23 ;
      RECT 5.875 0.66 5.965 1.23 ;
      RECT 5.44 0.66 5.53 1.065 ;
      RECT 6.235 0.675 6.94 0.765 ;
      RECT 4.745 0.66 5.965 0.75 ;
      RECT 5.625 0.325 5.715 0.75 ;
      RECT 4.325 0.25 4.415 0.965 ;
      RECT 4.325 0.25 5.114 0.34 ;
      RECT 4.325 0.25 5.194 0.279 ;
      RECT 5.156 0.17 5.56 0.26 ;
      RECT 5.076 0.231 5.56 0.26 ;
      RECT 5.114 0.191 5.156 0.319 ;
      RECT 4.12 1.14 4.595 1.23 ;
      RECT 4.505 0.45 4.595 1.23 ;
      RECT 1.965 1.14 2.5 1.23 ;
      RECT 2.93 1.075 3.42 1.165 ;
      RECT 3.33 1.06 4.21 1.15 ;
      RECT 2.41 1.06 3.02 1.15 ;
      RECT 1.965 0.48 2.055 1.23 ;
      RECT 4.505 0.93 5.325 1.02 ;
      RECT 4.505 0.45 5.405 0.54 ;
      RECT 5.265 0.35 5.405 0.54 ;
      RECT 3.33 0.88 4.03 0.97 ;
      RECT 3.94 0.29 4.03 0.97 ;
      RECT 2.355 0.25 2.445 0.635 ;
      RECT 3.37 0.29 4.18 0.38 ;
      RECT 4.03 0.17 4.18 0.38 ;
      RECT 2.355 0.25 3.01 0.34 ;
      RECT 3.37 0.17 3.46 0.38 ;
      RECT 2.92 0.17 3.46 0.26 ;
      RECT 3.125 0.35 3.215 0.985 ;
      RECT 3.76 0.47 3.85 0.655 ;
      RECT 3.125 0.47 3.85 0.56 ;
      RECT 3.1 0.35 3.24 0.55 ;
      RECT 2.56 0.46 3.24 0.55 ;
      RECT 2.175 0.325 2.265 0.985 ;
      RECT 2.175 0.74 2.815 0.83 ;
      RECT 2.725 0.685 3.02 0.775 ;
      RECT 0.695 1.06 1.87 1.15 ;
      RECT 1.78 0.17 1.87 1.15 ;
      RECT 1.78 0.17 1.925 0.37 ;
      RECT 0.88 0.25 1.46 0.34 ;
      RECT 0.545 0.22 1.015 0.335 ;
      RECT 1.37 0.17 1.925 0.26 ;
      RECT 0.87 0.88 1.69 0.97 ;
      RECT 1.6 0.35 1.69 0.97 ;
      RECT 0.87 0.725 0.96 0.97 ;
      RECT 0.43 0.725 0.96 0.815 ;
      RECT 0.43 0.48 0.52 0.815 ;
      RECT 1.55 0.35 1.69 0.44 ;
  END
END SDFFNX3H7R

MACRO SDFFQX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFQX0P5H7R 0 0 ;
  SIZE 6.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.4 1.48 ;
        RECT 5.845 1.015 5.935 1.48 ;
        RECT 4.7 1.225 4.84 1.48 ;
        RECT 3.46 1.225 3.6 1.48 ;
        RECT 2.63 1.225 2.77 1.48 ;
        RECT 1.19 1.21 1.33 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.4 0.08 ;
        RECT 5.845 -0.08 5.935 0.385 ;
        RECT 4.71 -0.08 4.85 0.295 ;
        RECT 3.56 -0.08 3.7 0.16 ;
        RECT 2.615 -0.08 2.755 0.16 ;
        RECT 1.075 -0.08 1.215 0.17 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.19 0.645 3.46 0.745 ;
      LAYER MET2 ;
        RECT 3.25 0.43 3.35 0.96 ;
      LAYER VIA1 ;
        RECT 3.255 0.655 3.345 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.025 0.31 6.185 1.03 ;
      LAYER MET2 ;
        RECT 6.05 0.43 6.15 0.96 ;
      LAYER VIA1 ;
        RECT 6.055 0.655 6.145 0.745 ;
    END
  END Q
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.33 0.455 1.42 0.625 ;
        RECT 0.64 0.455 1.42 0.545 ;
        RECT 0.64 0.455 0.73 0.605 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1 0.635 1.225 0.755 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.11 1.14 5.614 1.23 ;
      RECT 4.35 1.075 4.44 1.23 ;
      RECT 5.11 1.14 5.66 1.207 ;
      RECT 4.35 1.075 4.62 1.165 ;
      RECT 5.576 1.121 5.711 1.156 ;
      RECT 5.66 1.053 5.665 1.182 ;
      RECT 5.11 1.045 5.2 1.23 ;
      RECT 4.53 1.045 5.2 1.135 ;
      RECT 5.614 1.079 5.711 1.156 ;
      RECT 5.665 0.17 5.755 1.111 ;
      RECT 4.99 0.17 5.13 0.295 ;
      RECT 4.99 0.17 5.755 0.26 ;
      RECT 5.405 0.93 5.56 1.02 ;
      RECT 5.075 0.865 5.525 0.955 ;
      RECT 5.435 0.35 5.525 1.02 ;
      RECT 5.075 0.565 5.165 0.955 ;
      RECT 4.585 0.565 5.165 0.655 ;
      RECT 5.435 0.35 5.575 0.44 ;
      RECT 3.99 0.715 4.08 1.03 ;
      RECT 3.99 0.715 4.26 0.805 ;
      RECT 4.17 0.315 4.26 0.805 ;
      RECT 5.255 0.385 5.345 0.74 ;
      RECT 4.53 0.385 5.345 0.475 ;
      RECT 4.17 0.315 4.62 0.405 ;
      RECT 3.81 1.14 4.26 1.23 ;
      RECT 4.17 0.895 4.26 1.23 ;
      RECT 1.92 1.14 2.479 1.23 ;
      RECT 1.92 1.14 2.525 1.207 ;
      RECT 3.81 0.43 3.9 1.23 ;
      RECT 2.441 1.121 2.574 1.154 ;
      RECT 2.525 1.05 2.536 1.179 ;
      RECT 1.92 0.485 2.01 1.23 ;
      RECT 2.536 1.045 3.9 1.135 ;
      RECT 2.479 1.079 3.9 1.135 ;
      RECT 4.17 0.895 4.44 0.985 ;
      RECT 4.35 0.515 4.44 0.985 ;
      RECT 4.35 0.745 4.985 0.835 ;
      RECT 3.22 0.43 3.9 0.52 ;
      RECT 3.22 0.35 3.36 0.52 ;
      RECT 2.28 0.25 2.37 0.63 ;
      RECT 3.99 0.25 4.08 0.625 ;
      RECT 3.484 0.25 4.08 0.34 ;
      RECT 2.28 0.25 2.834 0.34 ;
      RECT 3.442 0.25 4.08 0.319 ;
      RECT 2.28 0.25 2.876 0.319 ;
      RECT 3.404 0.25 4.08 0.279 ;
      RECT 2.28 0.25 2.914 0.279 ;
      RECT 2.876 0.17 3.442 0.26 ;
      RECT 2.796 0.231 3.522 0.26 ;
      RECT 2.834 0.191 3.484 0.26 ;
      RECT 2.925 0.865 3.695 0.955 ;
      RECT 3.605 0.695 3.695 0.955 ;
      RECT 2.96 0.35 3.05 0.955 ;
      RECT 2.485 0.46 2.625 0.6 ;
      RECT 2.485 0.46 3.05 0.55 ;
      RECT 2.96 0.35 3.1 0.44 ;
      RECT 2.1 0.275 2.19 1.03 ;
      RECT 2.1 0.72 2.6 0.81 ;
      RECT 2.77 0.645 2.86 0.785 ;
      RECT 2.51 0.69 2.86 0.785 ;
      RECT 0.645 1.03 1.83 1.12 ;
      RECT 1.74 0.17 1.83 1.12 ;
      RECT 1.74 0.17 1.87 0.37 ;
      RECT 0.525 0.26 1.395 0.35 ;
      RECT 1.305 0.17 1.87 0.26 ;
      RECT 0.41 0.85 1.65 0.94 ;
      RECT 1.56 0.35 1.65 0.94 ;
      RECT 0.82 0.745 0.91 0.94 ;
      RECT 0.41 0.485 0.5 0.94 ;
      RECT 1.51 0.35 1.65 0.44 ;
  END
END SDFFQX0P5H7R

MACRO SDFFQX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFQX1H7R 0 0 ;
  SIZE 6.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.6 1.48 ;
        RECT 5.59 1.23 5.73 1.48 ;
        RECT 4.805 1.225 4.945 1.48 ;
        RECT 3.545 1.225 3.685 1.48 ;
        RECT 2.73 1.225 2.87 1.48 ;
        RECT 1.275 1.2 1.415 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.6 0.08 ;
        RECT 5.86 -0.08 6 0.16 ;
        RECT 5.005 -0.08 5.145 0.16 ;
        RECT 3.585 -0.08 3.725 0.16 ;
        RECT 2.715 -0.08 2.855 0.16 ;
        RECT 1.26 -0.08 1.4 0.17 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.35 0.625 3.575 0.745 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.055 0.345 6.29 0.435 ;
        RECT 5.95 0.695 6.145 0.785 ;
        RECT 6.055 0.345 6.145 0.785 ;
        RECT 5.95 0.695 6.04 0.985 ;
      LAYER MET2 ;
        RECT 6.05 0.23 6.15 0.76 ;
      LAYER VIA1 ;
        RECT 6.055 0.455 6.145 0.545 ;
    END
  END Q
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.036 0.645 1.52 0.735 ;
        RECT 0.93 0.626 1.074 0.652 ;
        RECT 0.93 0.6 1.036 0.652 ;
        RECT 1.022 0.645 1.52 0.728 ;
        RECT 0.884 0.57 1.022 0.606 ;
        RECT 0.976 0.645 1.52 0.698 ;
        RECT 0.884 0.524 0.976 0.606 ;
        RECT 0.625 0.478 0.93 0.545 ;
        RECT 0.625 0.455 0.884 0.545 ;
        RECT 0.846 0.524 0.976 0.564 ;
        RECT 0.625 0.455 0.73 0.605 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.115 0.455 1.385 0.555 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 4.415 1.045 4.555 1.23 ;
      RECT 4.415 1.045 5.86 1.135 ;
      RECT 5.77 0.269 5.86 1.135 ;
      RECT 2.38 0.25 2.47 0.575 ;
      RECT 4.931 0.255 5.435 0.345 ;
      RECT 3.504 0.25 3.879 0.34 ;
      RECT 2.38 0.25 2.944 0.34 ;
      RECT 5.764 0.198 5.77 0.326 ;
      RECT 4.885 0.193 4.931 0.321 ;
      RECT 3.462 0.25 3.921 0.319 ;
      RECT 2.38 0.25 2.986 0.319 ;
      RECT 5.726 0.269 5.86 0.304 ;
      RECT 5.345 0.195 5.764 0.285 ;
      RECT 4.847 0.17 4.885 0.279 ;
      RECT 3.424 0.25 3.959 0.279 ;
      RECT 2.38 0.25 3.024 0.279 ;
      RECT 5.77 0.224 5.816 1.135 ;
      RECT 3.921 0.17 4.885 0.26 ;
      RECT 4.931 0.236 4.97 0.345 ;
      RECT 3.879 0.191 3.921 0.319 ;
      RECT 2.906 0.231 3.542 0.26 ;
      RECT 3.841 0.231 4.932 0.26 ;
      RECT 4.931 0.216 4.932 0.345 ;
      RECT 2.944 0.191 3.504 0.26 ;
      RECT 2.986 0.17 3.462 0.26 ;
      RECT 4.525 0.865 5.68 0.955 ;
      RECT 5.59 0.375 5.68 0.955 ;
      RECT 4.525 0.72 4.665 0.955 ;
      RECT 5.525 0.375 5.68 0.465 ;
      RECT 4.055 0.35 4.145 1.03 ;
      RECT 5.285 0.605 5.5 0.75 ;
      RECT 5.285 0.45 5.375 0.75 ;
      RECT 4.871 0.45 5.375 0.54 ;
      RECT 4.855 0.404 4.871 0.532 ;
      RECT 4.809 0.373 4.855 0.501 ;
      RECT 4.771 0.431 4.909 0.459 ;
      RECT 4.055 0.35 4.809 0.44 ;
      RECT 3.85 1.14 4.325 1.23 ;
      RECT 4.235 0.53 4.325 1.23 ;
      RECT 2.02 1.14 2.579 1.23 ;
      RECT 2.02 1.14 2.625 1.207 ;
      RECT 2.986 1.115 3.36 1.205 ;
      RECT 2.954 1.061 2.986 1.189 ;
      RECT 2.916 1.115 3.36 1.154 ;
      RECT 3.85 0.43 3.94 1.23 ;
      RECT 2.541 1.121 2.674 1.154 ;
      RECT 2.625 1.05 2.636 1.179 ;
      RECT 2.02 0.485 2.11 1.23 ;
      RECT 3.27 1.045 3.94 1.135 ;
      RECT 2.636 1.045 2.954 1.135 ;
      RECT 2.579 1.096 3.024 1.135 ;
      RECT 2.579 1.079 2.986 1.135 ;
      RECT 4.794 0.63 5.14 0.72 ;
      RECT 4.778 0.584 4.794 0.712 ;
      RECT 4.732 0.553 4.778 0.681 ;
      RECT 4.694 0.611 4.832 0.639 ;
      RECT 4.235 0.53 4.732 0.62 ;
      RECT 3.295 0.43 3.94 0.52 ;
      RECT 3.295 0.35 3.385 0.52 ;
      RECT 3.065 0.35 3.155 1.025 ;
      RECT 3.065 0.835 3.76 0.925 ;
      RECT 3.67 0.675 3.76 0.925 ;
      RECT 2.585 0.46 3.155 0.55 ;
      RECT 2.2 0.24 2.29 1.03 ;
      RECT 2.2 0.725 2.965 0.815 ;
      RECT 0.525 1.02 1.93 1.11 ;
      RECT 1.84 0.17 1.93 1.11 ;
      RECT 0.525 0.26 1.479 0.35 ;
      RECT 1.84 0.17 1.97 0.345 ;
      RECT 0.525 0.26 1.525 0.327 ;
      RECT 0.525 0.26 1.569 0.279 ;
      RECT 1.531 0.17 1.97 0.26 ;
      RECT 1.441 0.241 1.97 0.26 ;
      RECT 1.525 0.173 1.531 0.301 ;
      RECT 1.479 0.199 1.97 0.26 ;
      RECT 0.41 0.84 1.7 0.93 ;
      RECT 1.61 0.35 1.7 0.93 ;
      RECT 0.825 0.795 0.965 0.93 ;
      RECT 0.41 0.485 0.5 0.93 ;
      RECT 1.61 0.35 1.75 0.44 ;
  END
END SDFFQX1H7R

MACRO SDFFQX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFQX2H7R 0 0 ;
  SIZE 6.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.6 1.48 ;
        RECT 6.17 1.035 6.26 1.48 ;
        RECT 5.605 1.23 5.745 1.48 ;
        RECT 4.805 1.225 4.945 1.48 ;
        RECT 3.545 1.225 3.685 1.48 ;
        RECT 2.73 1.225 2.87 1.48 ;
        RECT 1.25 1.21 1.39 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.6 0.08 ;
        RECT 6.36 -0.08 6.45 0.355 ;
        RECT 5.805 -0.08 5.945 0.16 ;
        RECT 4.955 -0.08 5.095 0.16 ;
        RECT 3.585 -0.08 3.725 0.16 ;
        RECT 2.715 -0.08 2.855 0.16 ;
        RECT 1.075 -0.08 1.215 0.17 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.35 0.635 3.575 0.755 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.91 0.455 6.2 0.545 ;
        RECT 6.11 0.235 6.2 0.545 ;
        RECT 5.91 0.455 6 1.11 ;
      LAYER MET2 ;
        RECT 6.05 0.23 6.15 0.76 ;
      LAYER VIA1 ;
        RECT 6.055 0.455 6.145 0.545 ;
    END
  END Q
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.036 0.645 1.52 0.735 ;
        RECT 0.93 0.626 1.074 0.652 ;
        RECT 0.93 0.6 1.036 0.652 ;
        RECT 1.022 0.645 1.52 0.728 ;
        RECT 0.884 0.57 1.022 0.606 ;
        RECT 0.976 0.645 1.52 0.698 ;
        RECT 0.884 0.524 0.976 0.606 ;
        RECT 0.625 0.478 0.93 0.545 ;
        RECT 0.625 0.455 0.884 0.545 ;
        RECT 0.846 0.524 0.976 0.564 ;
        RECT 0.625 0.455 0.73 0.605 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.115 0.455 1.385 0.555 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 4.415 1.045 4.555 1.215 ;
      RECT 4.415 1.045 5.81 1.135 ;
      RECT 5.72 0.274 5.81 1.135 ;
      RECT 2.38 0.25 2.47 0.58 ;
      RECT 4.881 0.255 5.385 0.345 ;
      RECT 3.504 0.25 3.879 0.34 ;
      RECT 2.38 0.25 2.934 0.34 ;
      RECT 5.709 0.2 5.72 0.329 ;
      RECT 4.835 0.193 4.881 0.321 ;
      RECT 3.462 0.25 3.921 0.319 ;
      RECT 2.38 0.25 2.976 0.319 ;
      RECT 5.671 0.274 5.81 0.304 ;
      RECT 5.295 0.195 5.709 0.285 ;
      RECT 4.797 0.17 4.835 0.279 ;
      RECT 3.424 0.25 3.959 0.279 ;
      RECT 2.38 0.25 3.014 0.279 ;
      RECT 5.72 0.229 5.766 1.135 ;
      RECT 3.921 0.17 4.835 0.26 ;
      RECT 4.881 0.236 4.92 0.345 ;
      RECT 3.879 0.191 3.921 0.319 ;
      RECT 2.896 0.231 3.542 0.26 ;
      RECT 3.841 0.231 4.882 0.26 ;
      RECT 4.881 0.216 4.882 0.345 ;
      RECT 2.934 0.191 3.504 0.26 ;
      RECT 2.976 0.17 3.462 0.26 ;
      RECT 4.59 0.865 5.63 0.955 ;
      RECT 5.54 0.375 5.63 0.955 ;
      RECT 4.59 0.79 4.68 0.955 ;
      RECT 5.49 0.375 5.63 0.465 ;
      RECT 4.055 0.35 4.145 1.03 ;
      RECT 5.36 0.584 5.45 0.75 ;
      RECT 5.325 0.498 5.36 0.627 ;
      RECT 5.279 0.458 5.325 0.586 ;
      RECT 5.279 0.539 5.406 0.586 ;
      RECT 5.241 0.435 5.279 0.544 ;
      RECT 4.805 0.435 5.279 0.525 ;
      RECT 4.759 0.373 4.805 0.501 ;
      RECT 4.721 0.35 4.759 0.459 ;
      RECT 4.055 0.35 4.759 0.44 ;
      RECT 4.055 0.416 4.844 0.44 ;
      RECT 4.055 0.396 4.806 0.44 ;
      RECT 3.85 1.14 4.325 1.23 ;
      RECT 4.235 0.53 4.325 1.23 ;
      RECT 2.02 1.14 2.579 1.23 ;
      RECT 2.02 1.14 2.625 1.207 ;
      RECT 2.946 1.075 3.36 1.165 ;
      RECT 2.916 1.075 3.36 1.15 ;
      RECT 3.85 0.43 3.94 1.23 ;
      RECT 2.541 1.121 2.674 1.154 ;
      RECT 2.625 1.05 2.636 1.179 ;
      RECT 2.02 0.485 2.11 1.23 ;
      RECT 3.27 1.045 3.94 1.135 ;
      RECT 2.579 1.079 3.94 1.135 ;
      RECT 2.636 1.045 2.954 1.135 ;
      RECT 2.625 1.06 2.984 1.135 ;
      RECT 4.728 0.615 5.14 0.705 ;
      RECT 4.682 0.553 4.728 0.681 ;
      RECT 4.644 0.615 5.14 0.639 ;
      RECT 4.235 0.53 4.682 0.62 ;
      RECT 4.235 0.596 4.767 0.62 ;
      RECT 4.235 0.576 4.729 0.62 ;
      RECT 3.295 0.43 3.94 0.52 ;
      RECT 3.295 0.35 3.385 0.52 ;
      RECT 3.065 0.35 3.155 0.985 ;
      RECT 3.065 0.865 3.76 0.955 ;
      RECT 3.67 0.635 3.76 0.955 ;
      RECT 2.585 0.46 3.155 0.55 ;
      RECT 2.2 0.24 2.29 1.035 ;
      RECT 2.2 0.685 2.965 0.775 ;
      RECT 0.525 1.03 1.93 1.12 ;
      RECT 1.84 0.17 1.93 1.12 ;
      RECT 0.525 0.26 1.479 0.35 ;
      RECT 1.84 0.17 1.97 0.345 ;
      RECT 0.525 0.26 1.525 0.327 ;
      RECT 0.525 0.26 1.569 0.279 ;
      RECT 1.531 0.17 1.97 0.26 ;
      RECT 1.441 0.241 1.97 0.26 ;
      RECT 1.525 0.173 1.531 0.301 ;
      RECT 1.479 0.199 1.97 0.26 ;
      RECT 0.41 0.84 1.7 0.93 ;
      RECT 1.61 0.35 1.7 0.93 ;
      RECT 0.825 0.795 0.965 0.93 ;
      RECT 0.41 0.485 0.5 0.93 ;
      RECT 1.61 0.35 1.75 0.44 ;
  END
END SDFFQX2H7R

MACRO SDFFQX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFQX3H7R 0 0 ;
  SIZE 7 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7 1.48 ;
        RECT 6.395 1.07 6.485 1.48 ;
        RECT 5.855 1.07 5.945 1.48 ;
        RECT 4.84 1.09 4.98 1.48 ;
        RECT 3.57 1.24 3.71 1.48 ;
        RECT 2.7 1.24 2.84 1.48 ;
        RECT 1.215 1.24 1.355 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7 0.08 ;
        RECT 6.395 -0.08 6.485 0.33 ;
        RECT 5.855 -0.08 5.945 0.33 ;
        RECT 4.85 -0.08 4.99 0.275 ;
        RECT 3.575 -0.08 3.715 0.16 ;
        RECT 2.645 -0.08 2.785 0.16 ;
        RECT 1.025 -0.08 1.165 0.16 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.255 0.625 3.475 0.775 ;
      LAYER MET2 ;
        RECT 3.25 0.43 3.35 0.96 ;
      LAYER VIA1 ;
        RECT 3.255 0.655 3.345 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.26 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.655 0.2 6.745 1.145 ;
        RECT 6.125 0.89 6.745 0.98 ;
        RECT 6.215 0.435 6.745 0.525 ;
        RECT 6.215 0.225 6.305 0.525 ;
        RECT 6.125 0.89 6.215 1.13 ;
        RECT 6.1 0.225 6.305 0.315 ;
      LAYER MET2 ;
        RECT 6.65 0.425 6.75 0.96 ;
      LAYER VIA1 ;
        RECT 6.655 0.655 6.745 0.745 ;
    END
  END Q
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.345 0.455 1.485 0.6 ;
        RECT 0.63 0.455 1.485 0.545 ;
        RECT 0.63 0.455 0.72 0.625 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.65 1.225 0.785 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.07 1.14 5.765 1.23 ;
      RECT 5.675 0.845 5.765 1.23 ;
      RECT 5.07 0.91 5.16 1.23 ;
      RECT 4.095 0.91 5.16 1 ;
      RECT 5.675 0.845 5.935 0.935 ;
      RECT 5.845 0.655 5.935 0.935 ;
      RECT 4.095 0.35 4.185 1 ;
      RECT 4.095 0.35 4.245 0.44 ;
      RECT 5.495 0.55 5.585 1.05 ;
      RECT 4.885 0.55 5.675 0.64 ;
      RECT 5.585 0.255 5.675 0.64 ;
      RECT 5.25 0.73 5.34 1.005 ;
      RECT 4.36 0.73 5.34 0.82 ;
      RECT 4.36 0.17 4.45 0.82 ;
      RECT 2.305 0.25 2.395 0.575 ;
      RECT 4.36 0.365 5.43 0.455 ;
      RECT 5.34 0.295 5.43 0.455 ;
      RECT 3.496 0.25 3.915 0.34 ;
      RECT 2.305 0.25 2.97 0.34 ;
      RECT 3.454 0.191 3.496 0.319 ;
      RECT 3.416 0.25 3.915 0.279 ;
      RECT 3.825 0.17 4.45 0.26 ;
      RECT 2.88 0.231 3.534 0.26 ;
      RECT 2.88 0.17 3.454 0.26 ;
      RECT 3.89 1.14 4.325 1.23 ;
      RECT 1.945 1.125 2.51 1.215 ;
      RECT 2.42 1.06 3.98 1.15 ;
      RECT 1.945 0.475 2.035 1.215 ;
      RECT 3.89 0.43 3.98 1.23 ;
      RECT 3.29 0.43 3.98 0.52 ;
      RECT 3.29 0.355 3.38 0.52 ;
      RECT 3.06 0.875 3.765 0.965 ;
      RECT 3.675 0.64 3.765 0.965 ;
      RECT 3.06 0.35 3.15 0.965 ;
      RECT 2.545 0.475 3.15 0.565 ;
      RECT 2.125 0.85 2.92 0.94 ;
      RECT 2.83 0.665 2.92 0.94 ;
      RECT 2.125 0.22 2.215 0.94 ;
      RECT 2.83 0.665 2.97 0.755 ;
      RECT 0.695 1.06 1.855 1.15 ;
      RECT 1.765 0.17 1.855 1.15 ;
      RECT 1.765 0.17 1.91 0.345 ;
      RECT 0.505 0.25 1.35 0.34 ;
      RECT 1.26 0.17 1.91 0.26 ;
      RECT 0.4 0.88 1.665 0.97 ;
      RECT 1.575 0.35 1.665 0.97 ;
      RECT 0.84 0.75 0.93 0.97 ;
      RECT 0.4 0.505 0.49 0.97 ;
  END
END SDFFQX3H7R

MACRO SDFFRQX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRQX0P5H7R 0 0 ;
  SIZE 6.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.4 1.48 ;
        RECT 5.99 1.07 6.08 1.48 ;
        RECT 5.245 1.05 5.335 1.48 ;
        RECT 3.755 1.185 3.845 1.48 ;
        RECT 3.26 1.005 3.35 1.48 ;
        RECT 2.11 1.195 2.2 1.48 ;
        RECT 1.215 1.095 1.355 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.4 0.08 ;
        RECT 5.99 -0.08 6.08 0.335 ;
        RECT 5.39 -0.08 5.48 0.345 ;
        RECT 3.235 -0.08 3.375 0.175 ;
        RECT 1.98 -0.08 2.07 0.33 ;
        RECT 1.125 -0.08 1.265 0.16 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.805 0.61 2.005 0.745 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.05 0.625 0.23 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.24 0.225 6.345 1.065 ;
      LAYER MET2 ;
        RECT 6.25 0.18 6.35 0.56 ;
      LAYER VIA1 ;
        RECT 6.255 0.255 6.345 0.345 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.2 0.845 5.47 0.945 ;
      LAYER MET2 ;
        RECT 5.25 0.625 5.35 1.16 ;
      LAYER VIA1 ;
        RECT 5.255 0.855 5.345 0.945 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.32 0.255 1.41 0.625 ;
        RECT 0.825 0.255 1.41 0.345 ;
        RECT 0.735 0.485 0.915 0.575 ;
        RECT 0.825 0.255 0.915 0.575 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.56 ;
      LAYER VIA1 ;
        RECT 0.855 0.255 0.945 0.345 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.455 1.225 0.59 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.74 0.925 5.9 1.065 ;
      RECT 5.81 0.44 5.9 1.065 ;
      RECT 4.99 0.44 5.9 0.53 ;
      RECT 5.74 0.295 5.83 0.53 ;
      RECT 5.47 1.045 5.65 1.135 ;
      RECT 5.56 0.63 5.65 1.135 ;
      RECT 4.705 0.35 4.795 1.045 ;
      RECT 4.705 0.63 5.72 0.72 ;
      RECT 4.57 0.35 4.795 0.44 ;
      RECT 3.755 0.17 3.845 0.365 ;
      RECT 5.14 0.17 5.23 0.35 ;
      RECT 3.755 0.17 5.23 0.26 ;
      RECT 4.525 1.135 5.005 1.225 ;
      RECT 4.915 0.81 5.005 1.225 ;
      RECT 4.525 0.594 4.615 1.225 ;
      RECT 4.115 0.96 4.615 1.05 ;
      RECT 2.55 0.96 3.05 1.05 ;
      RECT 2.96 0.825 3.05 1.05 ;
      RECT 4.115 0.825 4.205 1.05 ;
      RECT 2.55 0.17 2.64 1.05 ;
      RECT 2.96 0.825 4.205 0.915 ;
      RECT 4.51 0.518 4.525 0.647 ;
      RECT 4.464 0.488 4.51 0.616 ;
      RECT 4.464 0.549 4.571 0.616 ;
      RECT 4.426 0.549 4.571 0.574 ;
      RECT 4.24 0.465 4.464 0.555 ;
      RECT 2.97 0.285 3.64 0.375 ;
      RECT 2.97 0.17 3.06 0.375 ;
      RECT 2.55 0.17 3.06 0.26 ;
      RECT 4.295 0.78 4.435 0.87 ;
      RECT 4.295 0.645 4.385 0.87 ;
      RECT 4.06 0.645 4.385 0.735 ;
      RECT 4.06 0.35 4.15 0.735 ;
      RECT 3.12 0.465 4.15 0.555 ;
      RECT 4.01 0.35 4.15 0.555 ;
      RECT 3.935 1.14 4.345 1.23 ;
      RECT 3.44 1.14 3.585 1.23 ;
      RECT 3.495 1.005 3.585 1.23 ;
      RECT 3.935 1.005 4.025 1.23 ;
      RECT 3.495 1.005 4.025 1.095 ;
      RECT 2.73 0.645 2.87 0.87 ;
      RECT 2.73 0.645 3.955 0.735 ;
      RECT 2.73 0.35 2.82 0.87 ;
      RECT 2.73 0.35 2.87 0.44 ;
      RECT 2.32 1.14 2.975 1.23 ;
      RECT 1.685 1.14 2.02 1.23 ;
      RECT 1.93 1.015 2.02 1.23 ;
      RECT 2.32 0.42 2.41 1.23 ;
      RECT 1.93 1.015 2.41 1.105 ;
      RECT 1.73 0.42 2.41 0.51 ;
      RECT 1.73 0.25 1.82 0.51 ;
      RECT 1.441 0.96 1.84 1.05 ;
      RECT 1.75 0.835 1.84 1.05 ;
      RECT 1.434 0.918 1.441 1.047 ;
      RECT 0.32 0.935 1.104 1.025 ;
      RECT 1.396 0.96 1.84 1.024 ;
      RECT 0.32 0.935 1.124 1.015 ;
      RECT 1.086 0.915 1.434 1.005 ;
      RECT 0.32 0.941 1.479 1.005 ;
      RECT 1.066 0.925 1.441 1.005 ;
      RECT 0.32 0.295 0.41 1.025 ;
      RECT 1.75 0.835 2.195 0.925 ;
      RECT 2.105 0.695 2.195 0.925 ;
      RECT 0.32 0.295 0.715 0.385 ;
      RECT 1.52 0.735 1.66 0.87 ;
      RECT 0.885 0.735 1.025 0.835 ;
      RECT 0.5 0.735 1.66 0.825 ;
      RECT 1.5 0.275 1.59 0.825 ;
      RECT 0.5 0.5 0.59 0.825 ;
  END
END SDFFRQX0P5H7R

MACRO SDFFRQX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRQX1H7R 0 0 ;
  SIZE 6.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.6 1.48 ;
        RECT 6.06 1.04 6.15 1.48 ;
        RECT 5.29 1.05 5.38 1.48 ;
        RECT 3.74 1.21 3.88 1.48 ;
        RECT 3.305 1.055 3.395 1.48 ;
        RECT 2.165 1.195 2.255 1.48 ;
        RECT 1.235 1.095 1.375 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.6 0.08 ;
        RECT 5.94 -0.08 6.03 0.345 ;
        RECT 5.44 -0.08 5.53 0.345 ;
        RECT 3.28 -0.08 3.42 0.175 ;
        RECT 2.01 -0.08 2.1 0.33 ;
        RECT 1.135 -0.08 1.275 0.16 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.805 0.61 2.005 0.745 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.24 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.33 0.655 6.42 1.005 ;
        RECT 6.21 0.655 6.42 0.745 ;
        RECT 6.21 0.295 6.3 0.745 ;
      LAYER MET2 ;
        RECT 6.25 0.425 6.35 0.96 ;
      LAYER VIA1 ;
        RECT 6.255 0.655 6.345 0.745 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.225 0.845 5.505 0.945 ;
      LAYER MET2 ;
        RECT 5.25 0.625 5.35 1.16 ;
      LAYER VIA1 ;
        RECT 5.255 0.855 5.345 0.945 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.33 0.255 1.42 0.625 ;
        RECT 0.825 0.255 1.42 0.345 ;
        RECT 0.745 0.485 0.915 0.575 ;
        RECT 0.825 0.255 0.915 0.575 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.56 ;
      LAYER VIA1 ;
        RECT 0.855 0.255 0.945 0.345 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.445 1.225 0.58 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.785 0.93 5.96 1.02 ;
      RECT 5.87 0.44 5.96 1.02 ;
      RECT 5 0.44 5.96 0.53 ;
      RECT 5.67 0.295 5.76 0.53 ;
      RECT 5.535 1.03 5.685 1.12 ;
      RECT 5.595 0.62 5.685 1.12 ;
      RECT 4.74 0.35 4.83 1.05 ;
      RECT 4.74 0.62 5.78 0.71 ;
      RECT 4.58 0.35 4.83 0.44 ;
      RECT 3.81 0.17 3.9 0.375 ;
      RECT 5.105 0.17 5.195 0.35 ;
      RECT 3.81 0.17 5.195 0.26 ;
      RECT 4.56 1.14 5.04 1.23 ;
      RECT 4.95 0.81 5.04 1.23 ;
      RECT 4.56 0.639 4.65 1.23 ;
      RECT 4.15 0.96 4.65 1.05 ;
      RECT 2.595 0.96 3.135 1.05 ;
      RECT 3.045 0.85 3.135 1.05 ;
      RECT 4.15 0.85 4.24 1.05 ;
      RECT 2.595 0.17 2.685 1.05 ;
      RECT 3.045 0.85 4.24 0.94 ;
      RECT 4.525 0.553 4.56 0.682 ;
      RECT 4.479 0.513 4.525 0.641 ;
      RECT 4.479 0.594 4.606 0.641 ;
      RECT 4.441 0.49 4.479 0.599 ;
      RECT 4.335 0.49 4.479 0.58 ;
      RECT 3.07 0.285 3.67 0.375 ;
      RECT 3.58 0.23 3.67 0.375 ;
      RECT 3.07 0.17 3.16 0.375 ;
      RECT 2.595 0.17 3.16 0.26 ;
      RECT 4.33 0.78 4.47 0.87 ;
      RECT 4.319 0.675 4.33 0.804 ;
      RECT 4.319 0.749 4.42 0.804 ;
      RECT 4.281 0.749 4.42 0.779 ;
      RECT 4.13 0.67 4.319 0.76 ;
      RECT 4.13 0.704 4.376 0.76 ;
      RECT 4.13 0.35 4.22 0.76 ;
      RECT 3.165 0.465 4.22 0.555 ;
      RECT 4.075 0.35 4.22 0.555 ;
      RECT 3.97 1.14 4.375 1.23 ;
      RECT 3.51 1.14 3.65 1.23 ;
      RECT 3.56 1.03 3.65 1.23 ;
      RECT 3.97 1.03 4.06 1.23 ;
      RECT 3.56 1.03 4.06 1.12 ;
      RECT 2.775 0.645 2.915 0.87 ;
      RECT 2.775 0.645 4.035 0.735 ;
      RECT 2.775 0.35 2.865 0.87 ;
      RECT 2.775 0.35 2.915 0.44 ;
      RECT 2.365 1.14 3.02 1.23 ;
      RECT 1.695 1.14 2.075 1.23 ;
      RECT 1.985 1.015 2.075 1.23 ;
      RECT 2.365 0.42 2.455 1.23 ;
      RECT 1.985 1.015 2.455 1.105 ;
      RECT 1.74 0.42 2.455 0.51 ;
      RECT 1.74 0.255 1.83 0.51 ;
      RECT 0.33 0.965 1.099 1.055 ;
      RECT 1.461 0.96 1.895 1.05 ;
      RECT 1.805 0.835 1.895 1.05 ;
      RECT 1.454 0.918 1.461 1.047 ;
      RECT 1.416 0.96 1.895 1.024 ;
      RECT 0.33 0.965 1.149 1.024 ;
      RECT 1.111 0.915 1.454 1.005 ;
      RECT 1.099 0.921 1.111 1.049 ;
      RECT 0.33 0.275 0.42 1.055 ;
      RECT 1.061 0.946 1.499 1.005 ;
      RECT 1.461 0.941 1.499 1.05 ;
      RECT 1.805 0.835 2.225 0.925 ;
      RECT 2.135 0.665 2.225 0.925 ;
      RECT 0.33 0.275 0.725 0.365 ;
      RECT 1.575 0.735 1.715 0.87 ;
      RECT 0.895 0.735 1.035 0.835 ;
      RECT 0.51 0.735 1.715 0.825 ;
      RECT 1.51 0.275 1.6 0.825 ;
      RECT 0.51 0.5 0.6 0.825 ;
  END
END SDFFRQX1H7R

MACRO SDFFRQX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRQX2H7R 0 0 ;
  SIZE 6.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.6 1.48 ;
        RECT 6.14 1.06 6.23 1.48 ;
        RECT 5.38 1.035 5.47 1.48 ;
        RECT 3.92 1.21 4.06 1.48 ;
        RECT 3.355 1.185 3.445 1.48 ;
        RECT 2.07 1.195 2.16 1.48 ;
        RECT 1.235 1.095 1.375 1.48 ;
        RECT 0.07 1.005 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.6 0.08 ;
        RECT 6.41 -0.08 6.5 0.34 ;
        RECT 5.91 -0.08 6 0.34 ;
        RECT 5.43 -0.08 5.52 0.345 ;
        RECT 3.33 -0.08 3.47 0.175 ;
        RECT 2.01 -0.08 2.1 0.33 ;
        RECT 1.135 -0.08 1.275 0.16 ;
        RECT 0.07 -0.08 0.16 0.37 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.805 0.61 2.005 0.745 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.24 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.39 0.655 6.48 1.185 ;
        RECT 6.16 0.655 6.48 0.745 ;
        RECT 6.16 0.205 6.25 0.745 ;
      LAYER MET2 ;
        RECT 6.25 0.425 6.35 0.96 ;
      LAYER VIA1 ;
        RECT 6.255 0.655 6.345 0.745 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.405 0.81 5.605 0.945 ;
      LAYER MET2 ;
        RECT 5.45 0.625 5.55 1.16 ;
      LAYER VIA1 ;
        RECT 5.455 0.855 5.545 0.945 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.33 0.255 1.42 0.645 ;
        RECT 0.825 0.255 1.42 0.345 ;
        RECT 0.745 0.485 0.915 0.575 ;
        RECT 0.825 0.255 0.915 0.575 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.56 ;
      LAYER VIA1 ;
        RECT 0.855 0.255 0.945 0.345 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.455 1.225 0.59 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.88 0.925 6.035 1.065 ;
      RECT 5.945 0.44 6.035 1.065 ;
      RECT 5.025 0.44 6.035 0.53 ;
      RECT 5.66 0.25 5.75 0.53 ;
      RECT 5.625 1.04 5.785 1.13 ;
      RECT 5.695 0.62 5.785 1.13 ;
      RECT 4.81 0.35 4.9 1.05 ;
      RECT 4.81 0.62 5.855 0.71 ;
      RECT 4.635 0.35 4.9 0.44 ;
      RECT 3.91 0.17 4 0.375 ;
      RECT 5.16 0.17 5.25 0.345 ;
      RECT 3.91 0.17 5.25 0.26 ;
      RECT 4.6 1.14 5.13 1.23 ;
      RECT 5.04 0.81 5.13 1.23 ;
      RECT 4.6 0.53 4.69 1.23 ;
      RECT 4.291 0.96 4.69 1.05 ;
      RECT 2.645 0.96 3.044 1.05 ;
      RECT 4.286 0.919 4.291 1.048 ;
      RECT 2.645 0.96 3.09 1.027 ;
      RECT 4.24 0.894 4.286 1.022 ;
      RECT 4.194 0.848 4.24 0.976 ;
      RECT 4.194 0.941 4.329 0.976 ;
      RECT 3.006 0.941 3.136 0.981 ;
      RECT 2.645 0.17 2.735 1.05 ;
      RECT 3.044 0.899 3.141 0.956 ;
      RECT 4.156 0.825 4.194 0.934 ;
      RECT 3.044 0.899 3.179 0.934 ;
      RECT 3.141 0.825 4.194 0.915 ;
      RECT 3.136 0.827 3.141 0.956 ;
      RECT 3.09 0.853 4.24 0.915 ;
      RECT 4.455 0.53 4.69 0.62 ;
      RECT 3.12 0.285 3.77 0.375 ;
      RECT 3.68 0.23 3.77 0.375 ;
      RECT 3.12 0.17 3.21 0.375 ;
      RECT 2.645 0.17 3.21 0.26 ;
      RECT 4.37 0.755 4.51 0.87 ;
      RECT 4.365 0.663 4.37 0.792 ;
      RECT 4.321 0.733 4.459 0.767 ;
      RECT 4.321 0.689 4.416 0.767 ;
      RECT 4.275 0.35 4.365 0.722 ;
      RECT 3.215 0.465 4.365 0.555 ;
      RECT 4.225 0.35 4.365 0.555 ;
      RECT 4.211 1.14 4.51 1.23 ;
      RECT 2.415 1.14 3.144 1.23 ;
      RECT 1.7 1.14 1.899 1.23 ;
      RECT 4.185 1.089 4.211 1.217 ;
      RECT 2.415 1.14 3.19 1.207 ;
      RECT 1.7 1.14 1.945 1.207 ;
      RECT 4.139 1.053 4.185 1.181 ;
      RECT 4.139 1.121 4.249 1.181 ;
      RECT 3.106 1.121 3.236 1.161 ;
      RECT 2.415 0.42 2.505 1.23 ;
      RECT 1.861 1.121 1.986 1.164 ;
      RECT 4.101 1.03 4.139 1.139 ;
      RECT 3.144 1.079 3.241 1.136 ;
      RECT 1.899 1.079 2.024 1.124 ;
      RECT 1.945 1.035 1.986 1.164 ;
      RECT 3.69 1.03 4.139 1.12 ;
      RECT 3.144 1.079 3.279 1.114 ;
      RECT 1.986 1.015 2.505 1.105 ;
      RECT 3.241 1.005 3.78 1.095 ;
      RECT 3.236 1.007 3.241 1.136 ;
      RECT 3.19 1.033 4.139 1.095 ;
      RECT 1.74 0.42 2.505 0.51 ;
      RECT 1.74 0.225 1.83 0.51 ;
      RECT 2.825 0.35 2.965 0.87 ;
      RECT 2.825 0.645 4.185 0.735 ;
      RECT 0.33 1.04 1.024 1.13 ;
      RECT 0.33 1.04 1.07 1.107 ;
      RECT 1.461 0.96 1.814 1.05 ;
      RECT 1.454 0.918 1.461 1.047 ;
      RECT 0.986 1.021 1.111 1.064 ;
      RECT 0.33 0.275 0.42 1.13 ;
      RECT 1.454 0.96 1.86 1.027 ;
      RECT 1.416 0.96 1.86 1.024 ;
      RECT 1.024 0.979 1.149 1.024 ;
      RECT 1.07 0.935 1.111 1.064 ;
      RECT 1.111 0.915 1.454 1.005 ;
      RECT 1.776 0.941 1.901 0.984 ;
      RECT 1.07 0.941 1.499 1.005 ;
      RECT 1.814 0.899 1.939 0.944 ;
      RECT 1.86 0.855 1.901 0.984 ;
      RECT 2.135 0.6 2.225 0.925 ;
      RECT 1.901 0.835 2.225 0.925 ;
      RECT 0.33 0.275 0.735 0.365 ;
      RECT 1.575 0.735 1.715 0.87 ;
      RECT 0.895 0.735 1.035 0.835 ;
      RECT 0.51 0.735 1.715 0.825 ;
      RECT 1.51 0.235 1.6 0.825 ;
      RECT 0.51 0.5 0.6 0.825 ;
  END
END SDFFRQX2H7R

MACRO SDFFRX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRX0P5H7R 0 0 ;
  SIZE 7.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7.2 1.48 ;
        RECT 6.775 1.05 6.865 1.48 ;
        RECT 5.925 1.05 6.015 1.48 ;
        RECT 5.205 0.995 5.295 1.48 ;
        RECT 3.44 1.14 3.58 1.48 ;
        RECT 2 1.225 2.14 1.48 ;
        RECT 1.19 1.225 1.33 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7.2 0.08 ;
        RECT 6.775 -0.08 6.865 0.33 ;
        RECT 5.925 -0.08 6.015 0.35 ;
        RECT 5.01 -0.08 5.15 0.305 ;
        RECT 3.52 -0.08 3.66 0.185 ;
        RECT 1.975 -0.08 2.065 0.33 ;
        RECT 1.165 -0.08 1.255 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.885 0.455 2.175 0.555 ;
      LAYER MET2 ;
        RECT 2.05 0.23 2.15 0.76 ;
      LAYER VIA1 ;
        RECT 2.055 0.455 2.145 0.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.585 0.19 0.785 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.035 0.255 7.145 1.045 ;
      LAYER MET2 ;
        RECT 7.04 0.625 7.14 1.16 ;
      LAYER VIA1 ;
        RECT 7.045 0.855 7.135 0.945 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.285 0.255 6.375 1.045 ;
        RECT 6.18 0.255 6.375 0.345 ;
      LAYER MET2 ;
        RECT 6.25 0.18 6.35 0.56 ;
      LAYER VIA1 ;
        RECT 6.255 0.255 6.345 0.345 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.745 0.63 5.98 0.745 ;
      LAYER MET2 ;
        RECT 5.85 0.43 5.95 0.96 ;
      LAYER VIA1 ;
        RECT 5.855 0.655 5.945 0.745 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.33 0.425 1.42 0.605 ;
        RECT 0.855 0.425 1.42 0.515 ;
        RECT 0.695 0.49 0.945 0.58 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.625 1.235 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 6.105 1.14 6.615 1.23 ;
      RECT 6.525 0.295 6.615 1.23 ;
      RECT 5.385 1.135 5.835 1.225 ;
      RECT 5.745 0.87 5.835 1.225 ;
      RECT 6.105 0.87 6.195 1.23 ;
      RECT 5.385 0.76 5.475 1.225 ;
      RECT 5.745 0.87 6.195 0.96 ;
      RECT 4.835 0.76 5.475 0.85 ;
      RECT 6.525 0.705 6.945 0.795 ;
      RECT 6.855 0.655 6.945 0.795 ;
      RECT 4.4 0.78 4.54 0.87 ;
      RECT 4.4 0.215 4.49 0.87 ;
      RECT 6.075 0.445 6.165 0.68 ;
      RECT 5.745 0.445 6.165 0.535 ;
      RECT 4.83 0.395 5.375 0.485 ;
      RECT 5.285 0.17 5.375 0.485 ;
      RECT 5.745 0.17 5.835 0.535 ;
      RECT 4.83 0.215 4.92 0.485 ;
      RECT 4.4 0.215 4.92 0.305 ;
      RECT 5.285 0.17 5.835 0.26 ;
      RECT 5.565 0.35 5.655 1.045 ;
      RECT 5.13 0.58 5.655 0.67 ;
      RECT 5.515 0.35 5.655 0.44 ;
      RECT 3.67 1.14 5.045 1.23 ;
      RECT 4.955 0.96 5.045 1.23 ;
      RECT 2.77 1.14 3.23 1.23 ;
      RECT 3.14 0.96 3.23 1.23 ;
      RECT 2.77 0.755 2.86 1.23 ;
      RECT 3.14 0.96 4.74 1.05 ;
      RECT 4.65 0.395 4.74 1.05 ;
      RECT 4.21 0.7 4.3 1.05 ;
      RECT 2.73 0.465 2.82 0.845 ;
      RECT 4.22 0.17 4.31 0.58 ;
      RECT 3.12 0.285 3.21 0.555 ;
      RECT 3.12 0.285 3.89 0.375 ;
      RECT 3.8 0.17 3.89 0.375 ;
      RECT 3.8 0.17 4.31 0.26 ;
      RECT 3.98 0.78 4.12 0.87 ;
      RECT 3.98 0.35 4.07 0.87 ;
      RECT 3.325 0.49 4.07 0.58 ;
      RECT 3.98 0.35 4.12 0.44 ;
      RECT 2.95 0.6 3.04 1.045 ;
      RECT 2.95 0.675 3.89 0.765 ;
      RECT 2.94 0.22 3.03 0.69 ;
      RECT 0.28 1.045 2.68 1.135 ;
      RECT 2.55 0.97 2.68 1.135 ;
      RECT 0.28 0.295 0.37 1.135 ;
      RECT 2.55 0.255 2.64 1.135 ;
      RECT 0.28 0.295 0.665 0.385 ;
      RECT 2.32 0.865 2.46 0.955 ;
      RECT 2.37 0.255 2.46 0.955 ;
      RECT 2.255 0.255 2.46 0.345 ;
      RECT 1.7 0.865 2.23 0.955 ;
      RECT 2.14 0.695 2.23 0.955 ;
      RECT 1.7 0.255 1.79 0.955 ;
      RECT 0.87 0.865 1.6 0.955 ;
      RECT 1.51 0.245 1.6 0.955 ;
      RECT 0.87 0.745 0.96 0.955 ;
      RECT 0.46 0.745 0.96 0.835 ;
      RECT 0.46 0.505 0.55 0.835 ;
      RECT 1.405 0.245 1.6 0.335 ;
  END
END SDFFRX0P5H7R

MACRO SDFFRX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRX1H7R 0 0 ;
  SIZE 7.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7.2 1.48 ;
        RECT 6.78 1.07 6.87 1.48 ;
        RECT 5.96 1.05 6.05 1.48 ;
        RECT 5.23 0.995 5.32 1.48 ;
        RECT 3.44 1.14 3.58 1.48 ;
        RECT 1.98 1.225 2.12 1.48 ;
        RECT 1.19 1.225 1.33 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7.2 0.08 ;
        RECT 6.78 -0.08 6.87 0.33 ;
        RECT 5.96 -0.08 6.05 0.33 ;
        RECT 5.045 -0.08 5.185 0.305 ;
        RECT 3.57 -0.08 3.71 0.185 ;
        RECT 1.975 -0.08 2.065 0.33 ;
        RECT 1.18 -0.08 1.27 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.89 0.425 2.145 0.58 ;
      LAYER MET2 ;
        RECT 2.05 0.23 2.15 0.76 ;
      LAYER VIA1 ;
        RECT 2.055 0.455 2.145 0.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.585 0.19 0.785 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.005 0.89 7.145 0.98 ;
        RECT 7.055 0.32 7.145 0.98 ;
        RECT 7.005 0.32 7.145 0.41 ;
      LAYER MET2 ;
        RECT 7.05 0.63 7.15 1.16 ;
      LAYER VIA1 ;
        RECT 7.055 0.855 7.145 0.945 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.32 0.255 6.41 0.98 ;
        RECT 6.185 0.255 6.41 0.345 ;
      LAYER MET2 ;
        RECT 6.25 0.18 6.35 0.56 ;
      LAYER VIA1 ;
        RECT 6.255 0.255 6.345 0.345 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.78 0.625 5.96 0.775 ;
      LAYER MET2 ;
        RECT 5.85 0.43 5.95 0.96 ;
      LAYER VIA1 ;
        RECT 5.855 0.655 5.945 0.745 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.33 0.425 1.42 0.605 ;
        RECT 0.855 0.425 1.42 0.515 ;
        RECT 0.695 0.49 0.945 0.58 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.625 1.235 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.41 1.14 5.87 1.23 ;
      RECT 5.78 0.87 5.87 1.23 ;
      RECT 6.14 1.105 6.62 1.195 ;
      RECT 6.53 0.295 6.62 1.195 ;
      RECT 5.41 0.755 5.5 1.23 ;
      RECT 6.14 0.87 6.23 1.195 ;
      RECT 5.78 0.87 6.23 0.96 ;
      RECT 4.865 0.755 5.5 0.845 ;
      RECT 6.53 0.655 6.965 0.795 ;
      RECT 4.44 0.78 4.58 0.87 ;
      RECT 4.44 0.215 4.53 0.87 ;
      RECT 6.11 0.44 6.2 0.68 ;
      RECT 5.78 0.44 6.2 0.53 ;
      RECT 4.865 0.395 5.41 0.485 ;
      RECT 5.32 0.17 5.41 0.485 ;
      RECT 5.78 0.17 5.87 0.53 ;
      RECT 4.865 0.215 4.955 0.485 ;
      RECT 4.44 0.215 4.955 0.305 ;
      RECT 5.32 0.17 5.87 0.26 ;
      RECT 5.6 0.35 5.69 1.05 ;
      RECT 5.135 0.575 5.69 0.665 ;
      RECT 5.55 0.35 5.69 0.665 ;
      RECT 3.67 1.14 5.045 1.23 ;
      RECT 4.955 0.96 5.045 1.23 ;
      RECT 2.7 1.14 3.23 1.23 ;
      RECT 3.14 0.96 3.23 1.23 ;
      RECT 2.7 0.51 2.79 1.23 ;
      RECT 3.14 0.96 4.775 1.05 ;
      RECT 4.685 0.395 4.775 1.05 ;
      RECT 4.215 0.7 4.305 1.05 ;
      RECT 2.285 0.17 2.375 0.955 ;
      RECT 4.26 0.17 4.35 0.6 ;
      RECT 3.12 0.17 3.21 0.555 ;
      RECT 3.12 0.285 3.89 0.375 ;
      RECT 3.8 0.17 3.89 0.375 ;
      RECT 2.225 0.17 2.375 0.345 ;
      RECT 3.8 0.17 4.35 0.26 ;
      RECT 2.225 0.17 3.21 0.26 ;
      RECT 3.98 0.78 4.12 0.87 ;
      RECT 3.98 0.35 4.07 0.87 ;
      RECT 3.325 0.49 4.07 0.58 ;
      RECT 3.98 0.35 4.12 0.44 ;
      RECT 2.94 0.355 3.03 1.03 ;
      RECT 2.94 0.675 3.89 0.765 ;
      RECT 2.89 0.355 3.03 0.445 ;
      RECT 0.28 1.045 2.61 1.135 ;
      RECT 2.52 0.355 2.61 1.135 ;
      RECT 0.28 0.295 0.37 1.135 ;
      RECT 2.495 0.355 2.635 0.445 ;
      RECT 0.28 0.295 0.665 0.385 ;
      RECT 1.7 0.84 2.175 0.93 ;
      RECT 2.085 0.695 2.175 0.93 ;
      RECT 1.7 0.255 1.79 0.93 ;
      RECT 0.87 0.865 1.61 0.955 ;
      RECT 1.52 0.24 1.61 0.955 ;
      RECT 0.87 0.745 0.96 0.955 ;
      RECT 0.46 0.745 0.96 0.835 ;
      RECT 0.46 0.505 0.55 0.835 ;
      RECT 1.405 0.24 1.61 0.33 ;
  END
END SDFFRX1H7R

MACRO SDFFRX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRX2H7R 0 0 ;
  SIZE 7.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7.4 1.48 ;
        RECT 6.825 1.07 6.915 1.48 ;
        RECT 5.985 1.035 6.075 1.48 ;
        RECT 5.4 1.225 5.54 1.48 ;
        RECT 4.265 1.22 4.405 1.48 ;
        RECT 3.71 1.22 3.85 1.48 ;
        RECT 2.495 1.225 2.635 1.48 ;
        RECT 1.985 1.225 2.125 1.48 ;
        RECT 1.19 1.225 1.33 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7.4 0.08 ;
        RECT 7.215 -0.08 7.305 0.34 ;
        RECT 6.715 -0.08 6.805 0.33 ;
        RECT 6.235 -0.08 6.325 0.21 ;
        RECT 5.58 -0.08 5.67 0.33 ;
        RECT 3.66 -0.08 3.8 0.185 ;
        RECT 2.46 -0.08 2.6 0.185 ;
        RECT 1.99 -0.08 2.08 0.33 ;
        RECT 1.18 -0.08 1.27 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.88 0.455 2.175 0.545 ;
        RECT 1.88 0.455 1.97 0.645 ;
      LAYER MET2 ;
        RECT 2.05 0.23 2.15 0.76 ;
      LAYER VIA1 ;
        RECT 2.055 0.455 2.145 0.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.585 0.19 0.785 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.345 0.518 6.435 0.925 ;
        RECT 6.278 0.473 6.391 0.534 ;
        RECT 6.232 0.439 6.345 0.488 ;
        RECT 6.324 0.518 6.435 0.568 ;
        RECT 6.186 0.406 6.324 0.442 ;
        RECT 6.186 0.36 6.278 0.442 ;
        RECT 6.14 0.314 6.232 0.396 ;
        RECT 5.825 0.268 6.186 0.345 ;
        RECT 5.825 0.245 6.14 0.345 ;
        RECT 6.112 0.314 6.232 0.359 ;
      LAYER MET2 ;
        RECT 5.85 0.18 5.95 0.56 ;
      LAYER VIA1 ;
        RECT 5.855 0.255 5.945 0.345 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.055 0.805 7.165 1.155 ;
        RECT 7.035 0.235 7.125 0.87 ;
        RECT 6.94 0.235 7.125 0.325 ;
      LAYER MET2 ;
        RECT 7.05 0.63 7.15 1.16 ;
      LAYER VIA1 ;
        RECT 7.055 0.855 7.145 0.945 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.645 1.045 5.785 1.23 ;
        RECT 5.625 1.045 5.785 1.145 ;
        RECT 5.1 1.045 5.785 1.135 ;
        RECT 4.74 1.095 5.19 1.185 ;
        RECT 4.74 0.68 4.83 1.185 ;
        RECT 4.215 0.68 4.83 0.77 ;
        RECT 4.215 0.63 4.305 0.77 ;
      LAYER MET2 ;
        RECT 5.65 0.84 5.75 1.22 ;
      LAYER VIA1 ;
        RECT 5.655 1.055 5.745 1.145 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.33 0.425 1.42 0.705 ;
        RECT 0.855 0.425 1.42 0.515 ;
        RECT 0.695 0.485 0.945 0.575 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 0.625 1.23 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 6.165 1.015 6.69 1.105 ;
      RECT 6.525 0.32 6.615 1.105 ;
      RECT 6.165 0.624 6.255 1.105 ;
      RECT 5.41 0.445 5.5 0.775 ;
      RECT 6.146 0.546 6.165 0.675 ;
      RECT 6.1 0.514 6.146 0.642 ;
      RECT 6.525 0.54 6.94 0.63 ;
      RECT 6.1 0.579 6.211 0.642 ;
      RECT 6.054 0.468 6.1 0.596 ;
      RECT 6.016 0.445 6.054 0.554 ;
      RECT 5.41 0.445 6.054 0.535 ;
      RECT 6.44 0.32 6.615 0.41 ;
      RECT 4.92 0.865 5.01 1.005 ;
      RECT 4.92 0.865 5.915 0.955 ;
      RECT 5.825 0.625 5.915 0.955 ;
      RECT 5.23 0.235 5.32 0.955 ;
      RECT 5.825 0.625 5.965 0.715 ;
      RECT 4.695 0.235 5.32 0.325 ;
      RECT 2.29 0.28 2.38 0.955 ;
      RECT 5.05 0.465 5.14 0.775 ;
      RECT 3.34 0.17 3.43 0.585 ;
      RECT 4.44 0.465 5.14 0.555 ;
      RECT 4.44 0.17 4.53 0.555 ;
      RECT 3.34 0.285 3.98 0.375 ;
      RECT 3.89 0.17 3.98 0.375 ;
      RECT 2.215 0.28 2.8 0.37 ;
      RECT 2.71 0.17 2.8 0.37 ;
      RECT 3.89 0.17 4.53 0.26 ;
      RECT 2.71 0.17 3.43 0.26 ;
      RECT 4 0.86 4.65 0.95 ;
      RECT 4.035 0.49 4.125 0.95 ;
      RECT 3.545 0.49 4.125 0.58 ;
      RECT 4.041 0.467 4.171 0.511 ;
      RECT 4.087 0.425 4.181 0.483 ;
      RECT 4.087 0.425 4.219 0.459 ;
      RECT 4.181 0.35 4.325 0.44 ;
      RECT 4.125 0.383 4.325 0.44 ;
      RECT 4.171 0.355 4.181 0.483 ;
      RECT 4.505 1.14 4.645 1.23 ;
      RECT 2.93 1.14 3.59 1.23 ;
      RECT 3.5 1.04 3.59 1.23 ;
      RECT 4.505 1.04 4.595 1.23 ;
      RECT 2.93 0.46 3.02 1.23 ;
      RECT 3.5 1.04 4.595 1.13 ;
      RECT 2.47 0.46 2.56 0.665 ;
      RECT 2.47 0.46 3.02 0.55 ;
      RECT 3.26 0.675 3.35 1.03 ;
      RECT 3.11 0.675 3.945 0.765 ;
      RECT 3.11 0.355 3.2 0.765 ;
      RECT 3.11 0.355 3.25 0.445 ;
      RECT 0.28 1.045 2.79 1.135 ;
      RECT 2.7 0.655 2.79 1.135 ;
      RECT 0.28 0.295 0.37 1.135 ;
      RECT 0.28 0.295 0.645 0.385 ;
      RECT 1.7 0.855 2.2 0.945 ;
      RECT 2.11 0.635 2.2 0.945 ;
      RECT 1.7 0.295 1.79 0.945 ;
      RECT 0.87 0.865 1.6 0.955 ;
      RECT 1.51 0.245 1.6 0.955 ;
      RECT 0.87 0.745 0.96 0.955 ;
      RECT 0.46 0.745 0.96 0.835 ;
      RECT 0.46 0.505 0.55 0.835 ;
      RECT 1.405 0.245 1.6 0.335 ;
  END
END SDFFRX2H7R

MACRO SDFFRX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRX3H7R 0 0 ;
  SIZE 8.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 8.4 1.48 ;
        RECT 8.07 1.055 8.16 1.48 ;
        RECT 7.51 1.07 7.6 1.48 ;
        RECT 6.925 1.035 7.015 1.48 ;
        RECT 6.205 1.035 6.295 1.48 ;
        RECT 5.615 1.225 5.755 1.48 ;
        RECT 4.495 1.22 4.635 1.48 ;
        RECT 3.945 1.22 4.085 1.48 ;
        RECT 2.69 1.225 2.83 1.48 ;
        RECT 2.195 1.225 2.335 1.48 ;
        RECT 1.365 1.225 1.505 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 8.4 0.08 ;
        RECT 7.96 -0.08 8.05 0.34 ;
        RECT 7.42 -0.08 7.51 0.34 ;
        RECT 6.475 -0.08 6.565 0.2 ;
        RECT 5.765 -0.08 5.905 0.325 ;
        RECT 3.875 -0.08 4.015 0.185 ;
        RECT 2.675 -0.08 2.815 0.185 ;
        RECT 2.17 -0.08 2.26 0.35 ;
        RECT 1.335 -0.08 1.475 0.305 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 2.085 0.455 2.375 0.545 ;
        RECT 2.085 0.455 2.175 0.645 ;
      LAYER MET2 ;
        RECT 2.25 0.23 2.35 0.76 ;
      LAYER VIA1 ;
        RECT 2.255 0.455 2.345 0.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.24 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.43 0.655 6.88 0.745 ;
        RECT 6.79 0.21 6.88 0.745 ;
        RECT 6.565 0.655 6.655 0.925 ;
        RECT 6.43 0.418 6.52 0.745 ;
        RECT 6.361 0.373 6.476 0.432 ;
        RECT 6.315 0.338 6.43 0.386 ;
        RECT 6.407 0.418 6.52 0.467 ;
        RECT 6.277 0.304 6.407 0.344 ;
        RECT 6.12 0.258 6.361 0.325 ;
        RECT 6.12 0.235 6.315 0.325 ;
      LAYER MET2 ;
        RECT 6.65 0.425 6.75 0.96 ;
      LAYER VIA1 ;
        RECT 6.655 0.655 6.745 0.745 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.78 0.455 8.31 0.545 ;
        RECT 8.22 0.2 8.31 0.545 ;
        RECT 7.78 0.375 7.87 1.155 ;
        RECT 7.69 0.2 7.78 0.465 ;
      LAYER MET2 ;
        RECT 7.85 0.23 7.95 0.76 ;
      LAYER VIA1 ;
        RECT 7.855 0.455 7.945 0.545 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.845 1.045 5.985 1.23 ;
        RECT 5.825 1.045 5.985 1.145 ;
        RECT 5.365 1.045 5.985 1.135 ;
        RECT 4.97 1.12 5.455 1.21 ;
        RECT 4.97 0.759 5.06 1.21 ;
        RECT 4.435 0.714 5.016 0.77 ;
        RECT 4.435 0.685 4.97 0.77 ;
        RECT 4.959 0.759 5.06 0.814 ;
        RECT 4.435 0.68 4.959 0.77 ;
        RECT 4.921 0.759 5.06 0.789 ;
        RECT 4.435 0.615 4.55 0.77 ;
      LAYER MET2 ;
        RECT 5.85 0.84 5.95 1.22 ;
      LAYER VIA1 ;
        RECT 5.855 1.055 5.945 1.145 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.515 0.41 1.605 0.705 ;
        RECT 1.055 0.41 1.605 0.5 ;
        RECT 0.87 0.485 1.145 0.575 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.225 0.63 1.425 0.765 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 6.385 1.015 6.835 1.105 ;
      RECT 6.745 0.845 6.835 1.105 ;
      RECT 6.385 0.845 6.475 1.105 ;
      RECT 7.185 0.34 7.275 0.985 ;
      RECT 6.745 0.845 7.275 0.935 ;
      RECT 6.25 0.845 6.475 0.935 ;
      RECT 6.25 0.494 6.34 0.935 ;
      RECT 5.63 0.415 5.72 0.775 ;
      RECT 7.185 0.54 7.635 0.63 ;
      RECT 6.239 0.42 6.25 0.549 ;
      RECT 6.201 0.494 6.34 0.524 ;
      RECT 5.63 0.415 6.239 0.505 ;
      RECT 5.63 0.449 6.296 0.505 ;
      RECT 7.125 0.34 7.275 0.43 ;
      RECT 5.15 0.865 5.24 1.005 ;
      RECT 5.15 0.865 6.16 0.955 ;
      RECT 6.07 0.595 6.16 0.955 ;
      RECT 5.45 0.19 5.54 0.955 ;
      RECT 4.82 0.19 5.54 0.28 ;
      RECT 2.5 0.275 2.59 0.955 ;
      RECT 5.27 0.43 5.36 0.775 ;
      RECT 3.555 0.17 3.645 0.585 ;
      RECT 4.64 0.43 5.36 0.52 ;
      RECT 4.64 0.17 4.73 0.52 ;
      RECT 3.555 0.285 4.195 0.375 ;
      RECT 4.105 0.17 4.195 0.375 ;
      RECT 2.43 0.275 2.995 0.365 ;
      RECT 2.905 0.17 2.995 0.365 ;
      RECT 4.105 0.17 4.73 0.26 ;
      RECT 2.905 0.17 3.645 0.26 ;
      RECT 4.22 0.86 4.88 0.95 ;
      RECT 4.255 0.438 4.345 0.95 ;
      RECT 3.76 0.475 3.91 0.58 ;
      RECT 3.76 0.475 4.345 0.565 ;
      RECT 4.255 0.438 4.404 0.459 ;
      RECT 4.366 0.35 4.55 0.44 ;
      RECT 4.301 0.393 4.55 0.44 ;
      RECT 4.345 0.36 4.366 0.489 ;
      RECT 4.725 1.14 4.865 1.23 ;
      RECT 3.14 1.14 3.855 1.23 ;
      RECT 3.765 1.04 3.855 1.23 ;
      RECT 4.725 1.04 4.815 1.23 ;
      RECT 3.14 0.455 3.23 1.23 ;
      RECT 3.765 1.04 4.815 1.13 ;
      RECT 2.68 0.455 2.77 0.7 ;
      RECT 2.68 0.455 3.23 0.545 ;
      RECT 3.47 0.675 3.56 1.045 ;
      RECT 3.325 0.675 4.165 0.765 ;
      RECT 4.01 0.665 4.165 0.765 ;
      RECT 3.325 0.355 3.415 0.765 ;
      RECT 3.325 0.355 3.465 0.445 ;
      RECT 0.425 1.045 3 1.135 ;
      RECT 2.91 0.635 3 1.135 ;
      RECT 0.425 0.275 0.515 1.135 ;
      RECT 0.425 0.275 0.79 0.365 ;
      RECT 1.895 0.865 2.405 0.955 ;
      RECT 2.315 0.635 2.405 0.955 ;
      RECT 1.895 0.295 1.985 0.955 ;
      RECT 1.045 0.865 1.795 0.955 ;
      RECT 1.705 0.23 1.795 0.955 ;
      RECT 1.045 0.745 1.135 0.955 ;
      RECT 0.605 0.745 1.135 0.835 ;
      RECT 0.605 0.48 0.695 0.835 ;
      RECT 1.64 0.23 1.795 0.32 ;
  END
END SDFFRX3H7R

MACRO SDFFSQX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSQX1H7R 0 0 ;
  SIZE 7.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7.2 1.48 ;
        RECT 6.438 1.24 6.578 1.48 ;
        RECT 5.84 1.24 5.98 1.48 ;
        RECT 5.403 1.24 5.543 1.48 ;
        RECT 3.02 1.225 3.16 1.48 ;
        RECT 2.075 1.055 2.165 1.48 ;
        RECT 1.47 1.225 1.61 1.48 ;
        RECT 0.335 1.075 0.475 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7.2 0.08 ;
        RECT 6.661 -0.08 6.751 0.45 ;
        RECT 6.066 -0.08 6.206 0.16 ;
        RECT 5.16 -0.08 5.3 0.28 ;
        RECT 3.76 -0.08 3.85 0.345 ;
        RECT 3.02 -0.08 3.16 0.175 ;
        RECT 1.78 -0.08 1.92 0.32 ;
        RECT 1.28 -0.08 1.42 0.175 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.595 0.595 1.745 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.492 0.55 0.78 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.191 0.799 6.545 0.889 ;
        RECT 6.455 0.337 6.545 0.889 ;
        RECT 6.396 0.337 6.545 0.427 ;
        RECT 6.191 0.799 6.331 0.94 ;
      LAYER MET2 ;
        RECT 6.45 0.425 6.55 0.96 ;
      LAYER VIA1 ;
        RECT 6.455 0.655 6.545 0.745 ;
    END
  END Q
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.72 0.725 0.81 0.915 ;
        RECT 0.25 0.885 0.782 0.952 ;
        RECT 0.25 0.885 0.736 0.975 ;
        RECT 0.698 0.874 0.81 0.915 ;
        RECT 0.25 0.729 0.345 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.19 0.455 1.28 0.665 ;
        RECT 1.025 0.455 1.28 0.545 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END SI
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.855 0.57 5.975 0.795 ;
      LAYER MET2 ;
        RECT 5.85 0.43 5.95 0.96 ;
      LAYER VIA1 ;
        RECT 5.855 0.655 5.945 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 4.99 1.065 5.08 1.225 ;
      RECT 4.99 1.065 5.368 1.155 ;
      RECT 4.99 1.065 5.373 1.153 ;
      RECT 4.99 1.065 6.505 1.15 ;
      RECT 6.841 0.335 6.936 1.069 ;
      RECT 5.33 1.062 6.936 1.069 ;
      RECT 6.415 0.979 6.936 1.069 ;
      RECT 5.335 1.06 6.936 1.069 ;
      RECT 6.841 0.335 7.026 0.425 ;
      RECT 4.63 0.37 4.72 1.03 ;
      RECT 6.146 0.316 6.236 0.694 ;
      RECT 4.63 0.37 5.54 0.463 ;
      RECT 5.45 0.17 5.54 0.463 ;
      RECT 6.055 0.316 6.236 0.406 ;
      RECT 6.039 0.27 6.055 0.398 ;
      RECT 5.993 0.239 6.039 0.367 ;
      RECT 5.947 0.193 5.993 0.321 ;
      RECT 5.947 0.297 6.093 0.321 ;
      RECT 5.909 0.17 5.947 0.279 ;
      RECT 5.45 0.17 5.947 0.26 ;
      RECT 5.645 0.35 5.735 0.945 ;
      RECT 5.306 0.603 5.735 0.693 ;
      RECT 5.645 0.35 5.871 0.44 ;
      RECT 3.862 1.14 4.9 1.23 ;
      RECT 4.81 0.885 4.9 1.23 ;
      RECT 4.81 0.885 5.205 0.975 ;
      RECT 3.397 1.045 3.54 1.23 ;
      RECT 2.255 1.14 2.857 1.23 ;
      RECT 2.75 1.045 2.857 1.23 ;
      RECT 2.255 0.865 2.345 1.23 ;
      RECT 2.75 1.045 3.729 1.135 ;
      RECT 2.75 1.045 3.775 1.112 ;
      RECT 2.75 1.045 3.776 1.089 ;
      RECT 2.75 1.045 3.814 1.069 ;
      RECT 4.45 0.17 4.54 1.05 ;
      RECT 3.691 1.026 4.54 1.05 ;
      RECT 3.775 0.96 4.54 1.05 ;
      RECT 3.729 0.984 4.54 1.05 ;
      RECT 1.72 0.865 2.345 0.955 ;
      RECT 2.165 0.415 2.255 0.955 ;
      RECT 1.57 0.415 2.255 0.505 ;
      RECT 1.57 0.225 1.66 0.505 ;
      RECT 4.45 0.17 4.925 0.26 ;
      RECT 3.571 0.78 3.711 0.896 ;
      RECT 3.571 0.78 4.36 0.87 ;
      RECT 4.27 0.215 4.36 0.87 ;
      RECT 3.571 0.685 3.67 0.896 ;
      RECT 2.905 0.685 3.67 0.775 ;
      RECT 3.985 0.215 4.36 0.305 ;
      RECT 2.815 0.865 3.425 0.955 ;
      RECT 2.797 0.818 2.815 0.946 ;
      RECT 2.751 0.786 2.797 0.914 ;
      RECT 2.705 0.74 2.751 0.868 ;
      RECT 2.705 0.846 2.853 0.868 ;
      RECT 2.661 0.445 2.705 0.823 ;
      RECT 2.615 0.445 2.705 0.778 ;
      RECT 4.09 0.445 4.18 0.588 ;
      RECT 2.615 0.445 4.18 0.535 ;
      RECT 3.368 0.351 3.508 0.535 ;
      RECT 2.435 0.91 2.64 1.05 ;
      RECT 2.435 0.235 2.525 1.05 ;
      RECT 2.435 0.265 3.236 0.355 ;
      RECT 2.435 0.265 3.282 0.332 ;
      RECT 2.24 0.235 2.525 0.325 ;
      RECT 3.198 0.246 3.331 0.279 ;
      RECT 3.282 0.175 3.293 0.304 ;
      RECT 3.293 0.17 3.663 0.26 ;
      RECT 3.236 0.204 3.663 0.26 ;
      RECT 1.87 1.045 1.96 1.218 ;
      RECT 0.925 1.095 1.284 1.185 ;
      RECT 0.925 1.095 1.33 1.162 ;
      RECT 0.925 1.095 1.334 1.137 ;
      RECT 1.284 1.045 1.96 1.135 ;
      RECT 1.246 1.076 1.96 1.135 ;
      RECT 1.284 1.034 1.46 1.135 ;
      RECT 1.37 0.265 1.46 1.135 ;
      RECT 1.33 1.009 1.46 1.135 ;
      RECT 1.334 0.989 1.46 1.135 ;
      RECT 0.805 0.265 1.46 0.355 ;
      RECT 0.07 0.265 0.16 1.135 ;
      RECT 0.9 0.885 1.158 0.975 ;
      RECT 0.9 0.624 0.99 0.975 ;
      RECT 0.889 0.55 0.9 0.679 ;
      RECT 0.851 0.624 0.99 0.654 ;
      RECT 0.72 0.545 0.889 0.635 ;
      RECT 0.72 0.579 0.946 0.635 ;
      RECT 0.72 0.45 0.81 0.635 ;
      RECT 0.718 0.404 0.72 0.532 ;
      RECT 0.672 0.38 0.718 0.508 ;
      RECT 0.626 0.334 0.672 0.462 ;
      RECT 0.626 0.427 0.765 0.462 ;
      RECT 0.58 0.288 0.626 0.416 ;
      RECT 0.542 0.334 0.672 0.374 ;
      RECT 0.07 0.265 0.58 0.355 ;
  END
END SDFFSQX1H7R

MACRO SDFFSQX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSQX2H7R 0 0 ;
  SIZE 7.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7.2 1.48 ;
        RECT 6.438 1.24 6.578 1.48 ;
        RECT 5.84 1.24 5.98 1.48 ;
        RECT 5.375 1.24 5.515 1.48 ;
        RECT 3.025 1.225 3.165 1.48 ;
        RECT 2.075 1.055 2.165 1.48 ;
        RECT 1.47 1.225 1.61 1.48 ;
        RECT 0.31 1.225 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7.2 0.08 ;
        RECT 6.661 -0.08 6.751 0.45 ;
        RECT 6.066 -0.08 6.206 0.16 ;
        RECT 5.18 -0.08 5.32 0.175 ;
        RECT 3.765 -0.08 3.855 0.345 ;
        RECT 3.025 -0.08 3.165 0.175 ;
        RECT 1.78 -0.08 1.92 0.32 ;
        RECT 1.28 -0.08 1.42 0.175 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.595 0.595 1.745 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.492 0.55 0.78 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.191 0.799 6.545 0.889 ;
        RECT 6.455 0.337 6.545 0.889 ;
        RECT 6.396 0.337 6.545 0.427 ;
        RECT 6.191 0.799 6.331 0.94 ;
      LAYER MET2 ;
        RECT 6.45 0.425 6.55 0.96 ;
      LAYER VIA1 ;
        RECT 6.455 0.655 6.545 0.745 ;
    END
  END Q
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.883 0.82 0.985 ;
        RECT 0.73 0.73 0.82 0.985 ;
        RECT 0.25 0.73 0.345 0.985 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.19 0.455 1.28 0.635 ;
        RECT 1.025 0.455 1.28 0.545 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END SI
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.855 0.57 5.975 0.795 ;
      LAYER MET2 ;
        RECT 5.85 0.43 5.95 0.96 ;
      LAYER VIA1 ;
        RECT 5.855 0.655 5.945 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 5.01 1.065 5.1 1.225 ;
      RECT 5.01 1.065 5.318 1.155 ;
      RECT 5.01 1.065 5.323 1.153 ;
      RECT 5.01 1.065 6.505 1.15 ;
      RECT 6.841 0.335 6.936 1.069 ;
      RECT 5.28 1.062 6.936 1.069 ;
      RECT 6.415 0.979 6.936 1.069 ;
      RECT 5.285 1.06 6.936 1.069 ;
      RECT 6.841 0.335 7.026 0.425 ;
      RECT 4.65 0.37 4.74 1.025 ;
      RECT 6.146 0.316 6.236 0.694 ;
      RECT 4.65 0.37 5.56 0.463 ;
      RECT 5.47 0.17 5.56 0.463 ;
      RECT 6.055 0.316 6.236 0.406 ;
      RECT 6.039 0.27 6.055 0.398 ;
      RECT 5.993 0.239 6.039 0.367 ;
      RECT 5.947 0.193 5.993 0.321 ;
      RECT 5.947 0.297 6.093 0.321 ;
      RECT 5.909 0.17 5.947 0.279 ;
      RECT 5.47 0.17 5.947 0.26 ;
      RECT 5.645 0.553 5.74 0.945 ;
      RECT 5.65 0.35 5.74 0.945 ;
      RECT 5.275 0.553 5.74 0.643 ;
      RECT 5.65 0.35 5.871 0.44 ;
      RECT 3.862 1.14 4.92 1.23 ;
      RECT 4.83 0.885 4.92 1.23 ;
      RECT 4.83 0.885 5.225 0.975 ;
      RECT 3.397 1.045 3.54 1.23 ;
      RECT 2.255 1.14 2.857 1.23 ;
      RECT 2.75 1.045 2.857 1.23 ;
      RECT 2.255 0.865 2.345 1.23 ;
      RECT 2.75 1.045 3.729 1.135 ;
      RECT 2.75 1.045 3.775 1.112 ;
      RECT 2.75 1.045 3.776 1.089 ;
      RECT 2.75 1.045 3.814 1.069 ;
      RECT 4.47 0.17 4.56 1.05 ;
      RECT 3.691 1.026 4.56 1.05 ;
      RECT 3.775 0.96 4.56 1.05 ;
      RECT 3.729 0.984 4.56 1.05 ;
      RECT 1.72 0.865 2.345 0.955 ;
      RECT 2.165 0.415 2.255 0.955 ;
      RECT 1.57 0.415 2.255 0.505 ;
      RECT 1.57 0.225 1.66 0.505 ;
      RECT 4.47 0.17 4.945 0.26 ;
      RECT 3.571 0.685 3.711 0.896 ;
      RECT 3.571 0.78 4.38 0.87 ;
      RECT 4.29 0.24 4.38 0.87 ;
      RECT 2.91 0.685 3.711 0.775 ;
      RECT 3.99 0.24 4.38 0.33 ;
      RECT 2.83 0.865 3.43 0.955 ;
      RECT 2.797 0.81 2.83 0.939 ;
      RECT 2.751 0.771 2.797 0.899 ;
      RECT 2.751 0.846 2.868 0.899 ;
      RECT 2.705 0.725 2.751 0.853 ;
      RECT 2.661 0.445 2.705 0.808 ;
      RECT 2.615 0.445 2.705 0.763 ;
      RECT 4.11 0.445 4.2 0.588 ;
      RECT 2.615 0.445 4.2 0.535 ;
      RECT 3.373 0.351 3.513 0.535 ;
      RECT 2.435 0.91 2.64 1.05 ;
      RECT 2.435 0.235 2.525 1.05 ;
      RECT 2.435 0.265 3.241 0.355 ;
      RECT 2.435 0.265 3.287 0.332 ;
      RECT 2.26 0.235 2.525 0.325 ;
      RECT 3.203 0.246 3.336 0.279 ;
      RECT 3.287 0.175 3.298 0.304 ;
      RECT 3.298 0.17 3.67 0.26 ;
      RECT 3.241 0.204 3.67 0.26 ;
      RECT 1.87 1.045 1.96 1.218 ;
      RECT 0.829 1.076 1.373 1.166 ;
      RECT 0.829 1.076 1.404 1.151 ;
      RECT 1.37 1.045 1.96 1.135 ;
      RECT 1.335 1.058 1.96 1.135 ;
      RECT 1.37 0.265 1.46 1.135 ;
      RECT 0.805 0.265 1.46 0.355 ;
      RECT 0.07 0.265 0.16 1.056 ;
      RECT 0.93 0.895 1.158 0.985 ;
      RECT 0.93 0.65 1.02 0.985 ;
      RECT 0.898 0.566 0.93 0.694 ;
      RECT 0.86 0.605 0.976 0.659 ;
      RECT 0.72 0.55 0.898 0.64 ;
      RECT 0.72 0.45 0.81 0.64 ;
      RECT 0.718 0.404 0.72 0.532 ;
      RECT 0.672 0.38 0.718 0.508 ;
      RECT 0.626 0.334 0.672 0.462 ;
      RECT 0.626 0.427 0.765 0.462 ;
      RECT 0.58 0.288 0.626 0.416 ;
      RECT 0.542 0.334 0.672 0.374 ;
      RECT 0.07 0.265 0.58 0.355 ;
  END
END SDFFSQX2H7R

MACRO SDFFSQX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSQX3H7R 0 0 ;
  SIZE 7.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7.4 1.48 ;
        RECT 6.732 1.175 6.872 1.48 ;
        RECT 6.471 1.175 6.611 1.48 ;
        RECT 5.84 1.24 5.98 1.48 ;
        RECT 5.428 1.24 5.568 1.48 ;
        RECT 3.055 1.225 3.195 1.48 ;
        RECT 2.05 1.07 2.19 1.48 ;
        RECT 1.47 1.225 1.61 1.48 ;
        RECT 0.31 1.225 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7.4 0.08 ;
        RECT 6.894 -0.08 6.984 0.4 ;
        RECT 6.626 -0.08 6.766 0.16 ;
        RECT 6.066 -0.08 6.206 0.16 ;
        RECT 5.196 -0.08 5.336 0.28 ;
        RECT 3.796 -0.08 3.886 0.345 ;
        RECT 3.055 -0.08 3.195 0.175 ;
        RECT 1.78 -0.08 1.92 0.32 ;
        RECT 1.28 -0.08 1.42 0.175 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.595 0.595 1.745 0.775 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.492 0.55 0.78 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.191 0.799 6.745 0.905 ;
        RECT 6.655 0.337 6.745 0.905 ;
        RECT 6.346 0.337 6.745 0.427 ;
      LAYER MET2 ;
        RECT 6.65 0.425 6.75 0.96 ;
      LAYER VIA1 ;
        RECT 6.655 0.655 6.745 0.745 ;
    END
  END Q
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.72 0.73 0.81 0.95 ;
        RECT 0.25 0.933 0.766 0.995 ;
        RECT 0.677 0.914 0.81 0.95 ;
        RECT 0.715 0.892 0.72 1.021 ;
        RECT 0.25 0.933 0.715 1.023 ;
        RECT 0.25 0.73 0.345 1.023 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.19 0.455 1.28 0.595 ;
        RECT 1.025 0.455 1.28 0.545 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END SI
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.855 0.57 6.022 0.778 ;
      LAYER MET2 ;
        RECT 5.85 0.43 5.95 0.96 ;
      LAYER VIA1 ;
        RECT 5.855 0.655 5.945 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 5.063 1.075 5.153 1.225 ;
      RECT 5.063 1.075 5.358 1.165 ;
      RECT 5.063 1.075 5.36 1.164 ;
      RECT 5.063 1.075 5.398 1.144 ;
      RECT 7.074 0.335 7.169 1.085 ;
      RECT 5.32 1.056 7.169 1.085 ;
      RECT 5.875 0.995 7.169 1.085 ;
      RECT 5.358 1.036 7.169 1.085 ;
      RECT 5.36 1.035 5.965 1.125 ;
      RECT 7.074 0.335 7.259 0.425 ;
      RECT 4.666 0.37 4.756 1.019 ;
      RECT 6.121 0.579 6.461 0.669 ;
      RECT 6.121 0.316 6.236 0.669 ;
      RECT 4.666 0.37 5.576 0.463 ;
      RECT 5.486 0.17 5.576 0.463 ;
      RECT 6.055 0.316 6.236 0.406 ;
      RECT 6.039 0.27 6.055 0.398 ;
      RECT 5.993 0.239 6.039 0.367 ;
      RECT 5.947 0.193 5.993 0.321 ;
      RECT 5.947 0.297 6.093 0.321 ;
      RECT 5.909 0.17 5.947 0.279 ;
      RECT 5.486 0.17 5.947 0.26 ;
      RECT 5.645 0.553 5.765 0.945 ;
      RECT 5.675 0.35 5.765 0.945 ;
      RECT 5.31 0.553 5.765 0.643 ;
      RECT 5.675 0.35 5.871 0.44 ;
      RECT 3.862 1.14 4.973 1.23 ;
      RECT 4.883 0.885 4.973 1.23 ;
      RECT 4.883 0.885 5.288 0.975 ;
      RECT 3.397 1.045 3.54 1.23 ;
      RECT 2.322 1.14 2.857 1.23 ;
      RECT 2.75 1.045 2.857 1.23 ;
      RECT 2.322 0.865 2.412 1.23 ;
      RECT 2.75 1.045 3.729 1.135 ;
      RECT 2.75 1.045 3.775 1.112 ;
      RECT 2.75 1.045 3.776 1.089 ;
      RECT 2.75 1.045 3.814 1.069 ;
      RECT 4.486 0.17 4.576 1.05 ;
      RECT 3.691 1.026 4.576 1.05 ;
      RECT 3.775 0.96 4.576 1.05 ;
      RECT 3.729 0.984 4.576 1.05 ;
      RECT 1.72 0.865 2.412 0.955 ;
      RECT 2.193 0.415 2.283 0.955 ;
      RECT 1.57 0.415 2.283 0.505 ;
      RECT 1.57 0.225 1.66 0.505 ;
      RECT 4.486 0.17 4.64 0.26 ;
      RECT 3.571 0.78 3.711 0.896 ;
      RECT 3.571 0.78 4.396 0.87 ;
      RECT 4.306 0.215 4.396 0.87 ;
      RECT 3.571 0.685 3.67 0.896 ;
      RECT 2.965 0.685 3.67 0.775 ;
      RECT 2.965 0.625 3.055 0.775 ;
      RECT 4.033 0.215 4.396 0.305 ;
      RECT 2.86 0.865 3.466 0.955 ;
      RECT 2.818 0.806 2.86 0.934 ;
      RECT 2.772 0.762 2.818 0.89 ;
      RECT 2.772 0.846 2.898 0.89 ;
      RECT 2.728 0.445 2.772 0.845 ;
      RECT 2.682 0.445 2.772 0.8 ;
      RECT 4.126 0.445 4.216 0.605 ;
      RECT 2.682 0.445 4.216 0.535 ;
      RECT 3.403 0.351 3.543 0.535 ;
      RECT 2.502 0.91 2.66 1.05 ;
      RECT 2.502 0.235 2.592 1.05 ;
      RECT 2.855 0.265 3.271 0.355 ;
      RECT 2.855 0.265 3.317 0.332 ;
      RECT 2.25 0.235 2.945 0.325 ;
      RECT 3.233 0.246 3.366 0.279 ;
      RECT 3.317 0.175 3.328 0.304 ;
      RECT 3.328 0.17 3.706 0.26 ;
      RECT 3.271 0.204 3.706 0.26 ;
      RECT 1.87 1.045 1.96 1.218 ;
      RECT 0.909 1.09 1.289 1.18 ;
      RECT 0.909 1.09 1.334 1.158 ;
      RECT 1.289 1.045 1.96 1.135 ;
      RECT 1.251 1.071 1.96 1.135 ;
      RECT 1.289 1.029 1.46 1.135 ;
      RECT 1.37 0.265 1.46 1.135 ;
      RECT 1.334 0.989 1.46 1.135 ;
      RECT 0.805 0.265 1.46 0.355 ;
      RECT 0.07 0.265 0.16 1.071 ;
      RECT 1.01 0.728 1.1 1 ;
      RECT 0.993 0.651 1.01 0.79 ;
      RECT 0.947 0.62 0.993 0.758 ;
      RECT 0.947 0.683 1.056 0.758 ;
      RECT 0.901 0.574 0.947 0.712 ;
      RECT 0.855 0.528 0.901 0.666 ;
      RECT 0.853 0.445 0.855 0.642 ;
      RECT 0.807 0.574 0.947 0.618 ;
      RECT 0.72 0.445 0.855 0.595 ;
      RECT 0.677 0.378 0.72 0.512 ;
      RECT 0.631 0.334 0.677 0.467 ;
      RECT 0.631 0.422 0.765 0.467 ;
      RECT 0.585 0.288 0.631 0.421 ;
      RECT 0.542 0.334 0.677 0.377 ;
      RECT 0.07 0.265 0.585 0.355 ;
  END
END SDFFSQX3H7R

MACRO SDFFSRQX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRQX1H7R 0 0 ;
  SIZE 8.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 8.4 1.48 ;
        RECT 7.758 1.095 7.898 1.48 ;
        RECT 6.623 1.225 6.763 1.48 ;
        RECT 5.812 1.24 5.952 1.48 ;
        RECT 2.787 1.24 2.927 1.48 ;
        RECT 1.487 1.225 1.627 1.48 ;
        RECT 0.295 1.089 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 8.4 0.08 ;
        RECT 7.758 -0.08 7.898 0.305 ;
        RECT 6.948 -0.08 7.088 0.16 ;
        RECT 2.817 -0.08 2.957 0.28 ;
        RECT 1.258 -0.08 1.398 0.325 ;
        RECT 0.313 -0.08 0.453 0.175 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.223 0.45 3.442 0.62 ;
      LAYER MET2 ;
        RECT 3.25 0.23 3.35 0.76 ;
      LAYER VIA1 ;
        RECT 3.255 0.455 3.345 0.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.65 0.575 0.769 ;
        RECT 0.425 0.475 0.525 0.769 ;
        RECT 0.334 0.475 0.525 0.59 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 8.043 0.22 8.15 1.165 ;
      LAYER MET2 ;
        RECT 8.05 0.425 8.15 0.96 ;
      LAYER VIA1 ;
        RECT 8.055 0.655 8.145 0.745 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.399 0.569 6.624 0.768 ;
      LAYER MET2 ;
        RECT 6.45 0.425 6.55 0.96 ;
      LAYER VIA1 ;
        RECT 6.455 0.655 6.545 0.745 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.859 0.825 0.967 ;
        RECT 0.685 0.705 0.825 0.967 ;
        RECT 0.625 0.85 0.825 0.967 ;
        RECT 0.225 0.725 0.315 0.967 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.104 0.605 1.375 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END SI
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.023 0.45 7.248 0.661 ;
      LAYER MET2 ;
        RECT 7.05 0.23 7.15 0.76 ;
      LAYER VIA1 ;
        RECT 7.055 0.455 7.145 0.545 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 6.028 1.097 6.523 1.187 ;
      RECT 5.991 1.097 6.523 1.169 ;
      RECT 5.339 1.06 6.029 1.15 ;
      RECT 7.533 0.915 7.648 1.135 ;
      RECT 6.433 1.045 7.648 1.135 ;
      RECT 5.339 1.078 6.066 1.15 ;
      RECT 7.533 0.915 7.953 1.005 ;
      RECT 7.863 0.525 7.953 1.005 ;
      RECT 7.557 0.525 7.953 0.615 ;
      RECT 7.533 0.205 7.623 0.611 ;
      RECT 4.193 0.78 4.533 1.045 ;
      RECT 6.107 0.917 6.328 1.007 ;
      RECT 6.107 0.917 6.342 1 ;
      RECT 6.07 0.917 6.342 0.989 ;
      RECT 6.07 0.917 6.38 0.974 ;
      RECT 5.777 0.88 6.108 0.97 ;
      RECT 7.341 0.735 7.431 0.955 ;
      RECT 6.29 0.898 7.431 0.955 ;
      RECT 6.342 0.865 7.431 0.955 ;
      RECT 5.777 0.898 6.145 0.97 ;
      RECT 6.328 0.872 7.431 0.955 ;
      RECT 5.777 0.78 5.867 0.97 ;
      RECT 4.193 0.78 5.867 0.87 ;
      RECT 7.341 0.735 7.748 0.825 ;
      RECT 5.327 0.403 5.417 0.87 ;
      RECT 5.327 0.403 5.844 0.493 ;
      RECT 5.699 0.35 5.844 0.493 ;
      RECT 5.32 0.361 5.327 0.49 ;
      RECT 5.282 0.403 5.844 0.467 ;
      RECT 4.935 0.358 5.32 0.448 ;
      RECT 4.935 0.384 5.365 0.448 ;
      RECT 4.245 0.42 4.845 0.51 ;
      RECT 4.755 0.17 4.845 0.51 ;
      RECT 6.833 0.25 7.418 0.34 ;
      RECT 6.791 0.191 6.833 0.319 ;
      RECT 5.422 0.17 5.562 0.313 ;
      RECT 6.753 0.25 7.418 0.279 ;
      RECT 4.755 0.17 6.791 0.26 ;
      RECT 4.755 0.231 6.871 0.26 ;
      RECT 6.144 0.36 6.284 0.795 ;
      RECT 5.602 0.6 6.284 0.69 ;
      RECT 6.144 0.36 6.725 0.45 ;
      RECT 3.578 0.96 4.103 1.05 ;
      RECT 4.013 0.6 4.103 1.05 ;
      RECT 3.355 0.903 3.668 0.993 ;
      RECT 3.342 0.96 4.103 0.987 ;
      RECT 3.051 0.89 3.38 0.98 ;
      RECT 3.041 0.96 4.103 0.975 ;
      RECT 2.352 0.88 3.079 0.97 ;
      RECT 2.352 0.896 3.393 0.97 ;
      RECT 2.352 0.885 3.089 0.97 ;
      RECT 2.352 0.541 2.442 0.97 ;
      RECT 4.013 0.6 5.057 0.69 ;
      RECT 2.398 0.496 2.488 0.579 ;
      RECT 2.398 0.496 2.534 0.533 ;
      RECT 2.442 0.451 2.544 0.505 ;
      RECT 2.442 0.451 2.582 0.481 ;
      RECT 2.488 0.405 3.037 0.462 ;
      RECT 2.534 0.377 3.1 0.408 ;
      RECT 2.544 0.372 3.139 0.38 ;
      RECT 3.083 0.278 3.1 0.408 ;
      RECT 2.998 0.352 3.139 0.38 ;
      RECT 3.037 0.31 3.083 0.439 ;
      RECT 3.1 0.27 3.352 0.36 ;
      RECT 3.767 0.723 3.907 0.87 ;
      RECT 3.817 0.19 3.907 0.87 ;
      RECT 3.475 0.723 3.907 0.813 ;
      RECT 3.462 0.723 3.907 0.807 ;
      RECT 3.127 0.71 3.5 0.8 ;
      RECT 3.117 0.723 3.907 0.795 ;
      RECT 2.657 0.7 3.155 0.79 ;
      RECT 2.657 0.716 3.513 0.79 ;
      RECT 2.657 0.705 3.165 0.79 ;
      RECT 2.657 0.685 2.797 0.79 ;
      RECT 3.817 0.19 4.665 0.28 ;
      RECT 3.272 1.083 3.362 1.223 ;
      RECT 2.988 1.083 3.362 1.173 ;
      RECT 2.965 1.083 3.362 1.162 ;
      RECT 2.15 1.06 3.003 1.15 ;
      RECT 2.15 1.071 3.026 1.15 ;
      RECT 2.15 0.358 2.24 1.15 ;
      RECT 2.15 0.358 2.34 0.448 ;
      RECT 1.77 0.235 1.867 0.955 ;
      RECT 1.508 0.235 1.867 0.325 ;
      RECT 1.777 0.17 2.527 0.26 ;
      RECT 1.92 1.045 2.06 1.224 ;
      RECT 1.97 0.35 2.06 1.224 ;
      RECT 0.755 1.095 0.955 1.185 ;
      RECT 0.755 1.095 1.005 1.155 ;
      RECT 0.966 1.045 2.06 1.135 ;
      RECT 0.916 1.075 2.06 1.135 ;
      RECT 0.955 1.05 0.966 1.18 ;
      RECT 1.465 0.415 1.555 1.135 ;
      RECT 1.103 0.415 1.555 0.505 ;
      RECT 1.099 0.375 1.103 0.503 ;
      RECT 1.053 0.35 1.099 0.478 ;
      RECT 1.007 0.304 1.053 0.432 ;
      RECT 1.007 0.396 1.141 0.432 ;
      RECT 0.961 0.258 1.007 0.386 ;
      RECT 0.923 0.304 1.053 0.344 ;
      RECT 0.788 0.235 0.961 0.325 ;
      RECT 0.045 1.08 0.185 1.17 ;
      RECT 0.045 0.265 0.135 1.17 ;
      RECT 0.924 0.865 1.252 0.955 ;
      RECT 0.924 0.597 1.014 0.955 ;
      RECT 0.916 0.525 0.924 0.653 ;
      RECT 0.87 0.498 0.916 0.626 ;
      RECT 0.87 0.552 0.97 0.626 ;
      RECT 0.832 0.552 0.97 0.584 ;
      RECT 0.688 0.475 0.87 0.565 ;
      RECT 0.664 0.369 0.688 0.497 ;
      RECT 0.664 0.474 0.782 0.497 ;
      RECT 0.664 0.45 0.78 0.497 ;
      RECT 0.618 0.334 0.664 0.462 ;
      RECT 0.618 0.404 0.734 0.462 ;
      RECT 0.572 0.288 0.618 0.416 ;
      RECT 0.534 0.265 0.572 0.374 ;
      RECT 0.045 0.265 0.572 0.355 ;
      RECT 3.472 1.14 5.249 1.23 ;
  END
END SDFFSRQX1H7R

MACRO SDFFSRQX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRQX2H7R 0 0 ;
  SIZE 8.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 8.6 1.48 ;
        RECT 7.758 1.095 7.898 1.48 ;
        RECT 6.623 1.225 6.763 1.48 ;
        RECT 5.812 1.24 5.952 1.48 ;
        RECT 2.787 1.24 2.927 1.48 ;
        RECT 1.487 1.225 1.627 1.48 ;
        RECT 0.295 1.089 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 8.6 0.08 ;
        RECT 8.268 -0.08 8.408 0.32 ;
        RECT 7.758 -0.08 7.898 0.305 ;
        RECT 6.948 -0.08 7.088 0.16 ;
        RECT 2.817 -0.08 2.957 0.28 ;
        RECT 1.258 -0.08 1.398 0.325 ;
        RECT 0.313 -0.08 0.453 0.175 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.223 0.477 3.442 0.62 ;
        RECT 3.225 0.45 3.442 0.62 ;
      LAYER MET2 ;
        RECT 3.25 0.23 3.35 0.76 ;
      LAYER VIA1 ;
        RECT 3.255 0.455 3.345 0.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.65 0.575 0.769 ;
        RECT 0.425 0.475 0.525 0.769 ;
        RECT 0.334 0.475 0.525 0.59 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 8.043 0.22 8.15 1.165 ;
      LAYER MET2 ;
        RECT 8.05 0.425 8.15 0.96 ;
      LAYER VIA1 ;
        RECT 8.055 0.655 8.145 0.745 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.399 0.569 6.624 0.768 ;
      LAYER MET2 ;
        RECT 6.45 0.425 6.55 0.96 ;
      LAYER VIA1 ;
        RECT 6.455 0.655 6.545 0.745 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.859 0.825 0.967 ;
        RECT 0.685 0.705 0.825 0.967 ;
        RECT 0.625 0.85 0.825 0.967 ;
        RECT 0.225 0.725 0.315 0.967 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.104 0.605 1.375 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END SI
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.023 0.462 7.248 0.661 ;
        RECT 7.025 0.45 7.248 0.661 ;
      LAYER MET2 ;
        RECT 7.05 0.23 7.15 0.76 ;
      LAYER VIA1 ;
        RECT 7.055 0.455 7.145 0.545 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 6.028 1.097 6.523 1.187 ;
      RECT 5.991 1.097 6.523 1.169 ;
      RECT 5.339 1.06 6.029 1.15 ;
      RECT 7.533 0.915 7.623 1.135 ;
      RECT 6.433 1.045 7.623 1.135 ;
      RECT 5.339 1.078 6.066 1.15 ;
      RECT 7.533 0.915 7.953 1.005 ;
      RECT 7.863 0.525 7.953 1.005 ;
      RECT 7.533 0.525 7.953 0.615 ;
      RECT 7.533 0.209 7.623 0.615 ;
      RECT 4.193 0.78 4.533 1.045 ;
      RECT 6.107 0.917 6.328 1.007 ;
      RECT 6.107 0.917 6.342 1 ;
      RECT 6.07 0.917 6.342 0.989 ;
      RECT 6.07 0.917 6.38 0.974 ;
      RECT 5.777 0.88 6.108 0.97 ;
      RECT 7.341 0.735 7.431 0.955 ;
      RECT 6.29 0.898 7.431 0.955 ;
      RECT 6.342 0.865 7.431 0.955 ;
      RECT 5.777 0.898 6.145 0.97 ;
      RECT 6.328 0.872 7.431 0.955 ;
      RECT 5.777 0.78 5.867 0.97 ;
      RECT 4.193 0.78 5.867 0.87 ;
      RECT 7.341 0.735 7.748 0.825 ;
      RECT 5.327 0.403 5.417 0.87 ;
      RECT 5.327 0.403 5.844 0.493 ;
      RECT 5.699 0.35 5.844 0.493 ;
      RECT 5.32 0.361 5.327 0.49 ;
      RECT 5.282 0.403 5.844 0.467 ;
      RECT 4.935 0.358 5.32 0.448 ;
      RECT 4.935 0.384 5.365 0.448 ;
      RECT 4.245 0.42 4.845 0.51 ;
      RECT 4.755 0.17 4.845 0.51 ;
      RECT 6.833 0.25 7.418 0.34 ;
      RECT 6.791 0.191 6.833 0.319 ;
      RECT 5.422 0.17 5.562 0.313 ;
      RECT 6.753 0.25 7.418 0.279 ;
      RECT 4.755 0.17 6.791 0.26 ;
      RECT 4.755 0.231 6.871 0.26 ;
      RECT 6.144 0.36 6.284 0.795 ;
      RECT 5.602 0.6 6.284 0.69 ;
      RECT 6.144 0.36 6.725 0.45 ;
      RECT 3.578 0.96 4.103 1.05 ;
      RECT 4.013 0.6 4.103 1.05 ;
      RECT 3.355 0.903 3.668 0.993 ;
      RECT 3.342 0.96 4.103 0.987 ;
      RECT 3.051 0.89 3.38 0.98 ;
      RECT 3.041 0.96 4.103 0.975 ;
      RECT 2.352 0.88 3.079 0.97 ;
      RECT 2.352 0.896 3.393 0.97 ;
      RECT 2.352 0.885 3.089 0.97 ;
      RECT 2.352 0.541 2.442 0.97 ;
      RECT 4.013 0.6 5.057 0.69 ;
      RECT 2.398 0.496 2.488 0.579 ;
      RECT 2.398 0.496 2.534 0.533 ;
      RECT 2.442 0.451 2.544 0.505 ;
      RECT 2.442 0.451 2.582 0.481 ;
      RECT 2.488 0.405 3.037 0.462 ;
      RECT 2.534 0.377 3.1 0.408 ;
      RECT 2.544 0.372 3.139 0.38 ;
      RECT 3.083 0.278 3.1 0.408 ;
      RECT 2.998 0.352 3.139 0.38 ;
      RECT 3.037 0.31 3.083 0.439 ;
      RECT 3.1 0.27 3.352 0.36 ;
      RECT 3.767 0.723 3.907 0.87 ;
      RECT 3.817 0.19 3.907 0.87 ;
      RECT 3.475 0.723 3.907 0.813 ;
      RECT 3.462 0.723 3.907 0.807 ;
      RECT 3.127 0.71 3.5 0.8 ;
      RECT 3.117 0.723 3.907 0.795 ;
      RECT 2.657 0.7 3.155 0.79 ;
      RECT 2.657 0.716 3.513 0.79 ;
      RECT 2.657 0.705 3.165 0.79 ;
      RECT 2.657 0.685 2.797 0.79 ;
      RECT 3.817 0.19 4.665 0.28 ;
      RECT 3.272 1.083 3.362 1.223 ;
      RECT 2.988 1.083 3.362 1.173 ;
      RECT 2.965 1.083 3.362 1.162 ;
      RECT 2.15 1.06 3.003 1.15 ;
      RECT 2.15 1.071 3.026 1.15 ;
      RECT 2.15 0.358 2.24 1.15 ;
      RECT 2.15 0.358 2.34 0.448 ;
      RECT 1.77 0.235 1.867 0.955 ;
      RECT 1.508 0.235 1.867 0.325 ;
      RECT 1.777 0.17 2.527 0.26 ;
      RECT 1.92 1.045 2.06 1.224 ;
      RECT 1.97 0.35 2.06 1.224 ;
      RECT 0.755 1.095 0.955 1.185 ;
      RECT 0.755 1.095 1.005 1.155 ;
      RECT 0.966 1.045 2.06 1.135 ;
      RECT 0.916 1.075 2.06 1.135 ;
      RECT 0.955 1.05 0.966 1.18 ;
      RECT 1.465 0.415 1.555 1.135 ;
      RECT 1.103 0.415 1.555 0.505 ;
      RECT 1.099 0.375 1.103 0.503 ;
      RECT 1.053 0.35 1.099 0.478 ;
      RECT 1.007 0.304 1.053 0.432 ;
      RECT 1.007 0.396 1.141 0.432 ;
      RECT 0.961 0.258 1.007 0.386 ;
      RECT 0.923 0.304 1.053 0.344 ;
      RECT 0.788 0.235 0.961 0.325 ;
      RECT 0.045 1.08 0.185 1.17 ;
      RECT 0.045 0.265 0.135 1.17 ;
      RECT 0.924 0.865 1.252 0.955 ;
      RECT 0.924 0.597 1.014 0.955 ;
      RECT 0.916 0.525 0.924 0.653 ;
      RECT 0.87 0.498 0.916 0.626 ;
      RECT 0.87 0.552 0.97 0.626 ;
      RECT 0.832 0.552 0.97 0.584 ;
      RECT 0.688 0.475 0.87 0.565 ;
      RECT 0.664 0.369 0.688 0.497 ;
      RECT 0.664 0.474 0.782 0.497 ;
      RECT 0.664 0.45 0.78 0.497 ;
      RECT 0.618 0.334 0.664 0.462 ;
      RECT 0.618 0.404 0.734 0.462 ;
      RECT 0.572 0.288 0.618 0.416 ;
      RECT 0.534 0.265 0.572 0.374 ;
      RECT 0.045 0.265 0.572 0.355 ;
      RECT 3.472 1.14 5.249 1.23 ;
  END
END SDFFSRQX2H7R

MACRO SDFFSRQX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRQX3H7R 0 0 ;
  SIZE 8.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 8.6 1.48 ;
        RECT 8.268 1.08 8.408 1.48 ;
        RECT 7.758 1.095 7.898 1.48 ;
        RECT 6.623 1.225 6.763 1.48 ;
        RECT 5.812 1.24 5.952 1.48 ;
        RECT 2.787 1.24 2.927 1.48 ;
        RECT 1.487 1.225 1.627 1.48 ;
        RECT 0.295 1.089 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 8.6 0.08 ;
        RECT 8.268 -0.08 8.408 0.32 ;
        RECT 7.758 -0.08 7.898 0.305 ;
        RECT 6.948 -0.08 7.088 0.16 ;
        RECT 2.817 -0.08 2.957 0.28 ;
        RECT 1.258 -0.08 1.398 0.325 ;
        RECT 0.313 -0.08 0.453 0.175 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.223 0.477 3.442 0.62 ;
        RECT 3.225 0.45 3.442 0.62 ;
      LAYER MET2 ;
        RECT 3.25 0.23 3.35 0.76 ;
      LAYER VIA1 ;
        RECT 3.255 0.455 3.345 0.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.646 0.575 0.773 ;
        RECT 0.425 0.475 0.525 0.773 ;
        RECT 0.334 0.475 0.525 0.59 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 8.043 0.621 8.205 0.78 ;
        RECT 8.043 0.22 8.133 1.165 ;
      LAYER MET2 ;
        RECT 8.05 0.425 8.15 0.96 ;
      LAYER VIA1 ;
        RECT 8.055 0.655 8.145 0.745 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.399 0.569 6.624 0.768 ;
      LAYER MET2 ;
        RECT 6.45 0.425 6.55 0.96 ;
      LAYER VIA1 ;
        RECT 6.455 0.655 6.545 0.745 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.863 0.825 0.971 ;
        RECT 0.685 0.705 0.825 0.971 ;
        RECT 0.625 0.85 0.825 0.971 ;
        RECT 0.225 0.725 0.315 0.971 ;
      LAYER MET2 ;
        RECT 0.65 0.625 0.75 1.16 ;
      LAYER VIA1 ;
        RECT 0.655 0.855 0.745 0.945 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.104 0.605 1.375 0.775 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END SI
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.023 0.45 7.248 0.661 ;
      LAYER MET2 ;
        RECT 7.05 0.23 7.15 0.76 ;
      LAYER VIA1 ;
        RECT 7.055 0.455 7.145 0.545 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 6.028 1.097 6.523 1.187 ;
      RECT 5.991 1.097 6.523 1.169 ;
      RECT 5.339 1.06 6.029 1.15 ;
      RECT 7.533 0.915 7.623 1.135 ;
      RECT 6.433 1.045 7.623 1.135 ;
      RECT 5.339 1.078 6.066 1.15 ;
      RECT 7.533 0.915 7.953 1.005 ;
      RECT 7.863 0.525 7.953 1.005 ;
      RECT 7.533 0.525 7.953 0.615 ;
      RECT 7.533 0.209 7.623 0.615 ;
      RECT 4.193 0.78 4.533 1.045 ;
      RECT 6.107 0.917 6.328 1.007 ;
      RECT 6.107 0.917 6.342 1 ;
      RECT 6.07 0.917 6.342 0.989 ;
      RECT 6.07 0.917 6.38 0.974 ;
      RECT 5.777 0.88 6.108 0.97 ;
      RECT 7.341 0.735 7.431 0.955 ;
      RECT 6.29 0.898 7.431 0.955 ;
      RECT 6.342 0.865 7.431 0.955 ;
      RECT 5.777 0.898 6.145 0.97 ;
      RECT 6.328 0.872 7.431 0.955 ;
      RECT 5.777 0.78 5.867 0.97 ;
      RECT 4.193 0.78 5.867 0.87 ;
      RECT 7.341 0.735 7.748 0.825 ;
      RECT 5.327 0.403 5.417 0.87 ;
      RECT 5.327 0.403 5.844 0.493 ;
      RECT 5.699 0.35 5.844 0.493 ;
      RECT 5.32 0.361 5.327 0.49 ;
      RECT 5.282 0.403 5.844 0.467 ;
      RECT 4.935 0.358 5.32 0.448 ;
      RECT 4.935 0.384 5.365 0.448 ;
      RECT 4.245 0.42 4.845 0.51 ;
      RECT 4.755 0.17 4.845 0.51 ;
      RECT 6.833 0.25 7.418 0.34 ;
      RECT 6.791 0.191 6.833 0.319 ;
      RECT 5.422 0.17 5.562 0.313 ;
      RECT 6.753 0.25 7.418 0.279 ;
      RECT 4.755 0.17 6.791 0.26 ;
      RECT 4.755 0.231 6.871 0.26 ;
      RECT 6.144 0.36 6.284 0.795 ;
      RECT 5.602 0.6 6.284 0.69 ;
      RECT 6.144 0.36 6.725 0.45 ;
      RECT 3.578 0.96 4.103 1.05 ;
      RECT 4.013 0.6 4.103 1.05 ;
      RECT 3.355 0.903 3.668 0.993 ;
      RECT 3.342 0.96 4.103 0.987 ;
      RECT 3.051 0.89 3.38 0.98 ;
      RECT 3.041 0.96 4.103 0.975 ;
      RECT 2.352 0.88 3.079 0.97 ;
      RECT 2.352 0.896 3.393 0.97 ;
      RECT 2.352 0.885 3.089 0.97 ;
      RECT 2.352 0.541 2.442 0.97 ;
      RECT 4.013 0.6 5.057 0.69 ;
      RECT 2.398 0.496 2.488 0.579 ;
      RECT 2.398 0.496 2.534 0.533 ;
      RECT 2.442 0.451 2.544 0.505 ;
      RECT 2.442 0.451 2.582 0.481 ;
      RECT 2.488 0.405 3.037 0.462 ;
      RECT 2.534 0.377 3.1 0.408 ;
      RECT 2.544 0.372 3.139 0.38 ;
      RECT 3.083 0.278 3.1 0.408 ;
      RECT 2.998 0.352 3.139 0.38 ;
      RECT 3.037 0.31 3.083 0.439 ;
      RECT 3.1 0.27 3.352 0.36 ;
      RECT 3.767 0.723 3.907 0.87 ;
      RECT 3.817 0.19 3.907 0.87 ;
      RECT 3.475 0.723 3.907 0.813 ;
      RECT 3.462 0.723 3.907 0.807 ;
      RECT 3.127 0.71 3.5 0.8 ;
      RECT 3.117 0.723 3.907 0.795 ;
      RECT 2.657 0.7 3.155 0.79 ;
      RECT 2.657 0.716 3.513 0.79 ;
      RECT 2.657 0.705 3.165 0.79 ;
      RECT 2.657 0.685 2.797 0.79 ;
      RECT 3.817 0.19 4.665 0.28 ;
      RECT 3.272 1.083 3.362 1.223 ;
      RECT 2.988 1.083 3.362 1.173 ;
      RECT 2.965 1.083 3.362 1.162 ;
      RECT 2.15 1.06 3.003 1.15 ;
      RECT 2.15 1.071 3.026 1.15 ;
      RECT 2.15 0.358 2.24 1.15 ;
      RECT 2.15 0.358 2.34 0.448 ;
      RECT 1.77 0.235 1.867 0.955 ;
      RECT 1.508 0.235 1.867 0.325 ;
      RECT 1.777 0.17 2.527 0.26 ;
      RECT 1.92 1.045 2.06 1.224 ;
      RECT 1.97 0.35 2.06 1.224 ;
      RECT 0.755 1.095 0.955 1.185 ;
      RECT 0.755 1.095 1.005 1.155 ;
      RECT 0.966 1.045 2.06 1.135 ;
      RECT 0.916 1.075 2.06 1.135 ;
      RECT 0.955 1.05 0.966 1.18 ;
      RECT 1.465 0.415 1.555 1.135 ;
      RECT 1.103 0.415 1.555 0.505 ;
      RECT 1.099 0.375 1.103 0.503 ;
      RECT 1.053 0.35 1.099 0.478 ;
      RECT 1.007 0.304 1.053 0.432 ;
      RECT 1.007 0.396 1.141 0.432 ;
      RECT 0.961 0.258 1.007 0.386 ;
      RECT 0.923 0.304 1.053 0.344 ;
      RECT 0.788 0.235 0.961 0.325 ;
      RECT 0.045 1.08 0.185 1.17 ;
      RECT 0.045 0.265 0.135 1.17 ;
      RECT 0.924 0.865 1.252 0.955 ;
      RECT 0.924 0.597 1.014 0.955 ;
      RECT 0.916 0.525 0.924 0.653 ;
      RECT 0.87 0.498 0.916 0.626 ;
      RECT 0.87 0.552 0.97 0.626 ;
      RECT 0.832 0.552 0.97 0.584 ;
      RECT 0.688 0.475 0.87 0.565 ;
      RECT 0.664 0.369 0.688 0.497 ;
      RECT 0.664 0.474 0.782 0.497 ;
      RECT 0.664 0.45 0.78 0.497 ;
      RECT 0.618 0.334 0.664 0.462 ;
      RECT 0.618 0.404 0.734 0.462 ;
      RECT 0.572 0.288 0.618 0.416 ;
      RECT 0.534 0.265 0.572 0.374 ;
      RECT 0.045 0.265 0.572 0.355 ;
      RECT 3.472 1.14 5.249 1.23 ;
  END
END SDFFSRQX3H7R

MACRO SDFFSRX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRX0P5H7R 0 0 ;
  SIZE 8.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 8.8 1.48 ;
        RECT 8.065 1.028 8.155 1.48 ;
        RECT 7.35 1.24 7.49 1.48 ;
        RECT 6.386 1.24 6.526 1.48 ;
        RECT 5.385 1.24 5.525 1.48 ;
        RECT 2.807 1.24 2.947 1.48 ;
        RECT 1.466 1.225 1.606 1.48 ;
        RECT 0.381 1.095 0.521 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 8.8 0.08 ;
        RECT 8.065 -0.08 8.155 0.41 ;
        RECT 7.27 -0.08 7.41 0.305 ;
        RECT 6.103 -0.08 6.243 0.16 ;
        RECT 2.86 -0.08 3 0.16 ;
        RECT 1.378 -0.08 1.518 0.16 ;
        RECT 0.378 -0.08 0.518 0.305 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.728 0.625 1.95 0.775 ;
        RECT 1.728 0.59 1.945 0.795 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.622 0.631 0.808 ;
        RECT 0.43 0.622 0.631 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 8.315 0.63 8.575 0.75 ;
        RECT 8.315 0.286 8.405 1.082 ;
      LAYER MET2 ;
        RECT 8.45 0.43 8.55 0.96 ;
      LAYER VIA1 ;
        RECT 8.455 0.655 8.545 0.745 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.705 0.225 7.95 0.375 ;
        RECT 7.705 0.225 7.795 0.945 ;
      LAYER MET2 ;
        RECT 7.85 0.18 7.95 0.56 ;
      LAYER VIA1 ;
        RECT 7.855 0.255 7.945 0.345 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.225 0.45 6.375 0.55 ;
        RECT 6.205 0.455 6.295 0.749 ;
      LAYER MET2 ;
        RECT 6.25 0.225 6.35 0.76 ;
      LAYER VIA1 ;
        RECT 6.255 0.455 6.345 0.545 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.9 0.856 0.99 ;
        RECT 0.766 0.74 0.856 0.99 ;
        RECT 0.225 0.85 0.375 0.99 ;
        RECT 0.225 0.655 0.34 0.99 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.16 0.445 1.442 0.602 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END SI
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.465 0.45 6.775 0.628 ;
      LAYER MET2 ;
        RECT 6.65 0.225 6.75 0.76 ;
      LAYER VIA1 ;
        RECT 6.655 0.455 6.745 0.545 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 5.615 1.14 6.267 1.23 ;
      RECT 4.952 1.071 5.092 1.229 ;
      RECT 5.615 1.14 6.308 1.21 ;
      RECT 5.615 1.14 6.347 1.17 ;
      RECT 4.952 1.071 5.335 1.161 ;
      RECT 7.885 0.546 7.975 1.15 ;
      RECT 5.29 1.059 5.705 1.149 ;
      RECT 6.228 1.12 7.975 1.15 ;
      RECT 7.525 1.059 7.975 1.15 ;
      RECT 6.267 1.08 7.975 1.15 ;
      RECT 6.308 1.06 7.975 1.15 ;
      RECT 7.525 0.395 7.615 1.15 ;
      RECT 7.885 0.546 8.176 0.636 ;
      RECT 7.02 0.395 7.615 0.485 ;
      RECT 7.02 0.264 7.16 0.485 ;
      RECT 5.795 0.959 6.191 1.049 ;
      RECT 5.795 0.959 6.232 1.029 ;
      RECT 4.592 0.711 4.682 0.997 ;
      RECT 5.795 0.959 6.27 0.989 ;
      RECT 6.865 0.575 6.955 0.97 ;
      RECT 6.153 0.94 6.955 0.97 ;
      RECT 6.232 0.88 6.955 0.97 ;
      RECT 5.795 0.711 5.885 1.049 ;
      RECT 6.191 0.9 6.955 0.97 ;
      RECT 4.592 0.711 5.885 0.801 ;
      RECT 6.865 0.575 7.247 0.715 ;
      RECT 4.999 0.351 5.089 0.801 ;
      RECT 4.513 0.351 5.623 0.441 ;
      RECT 6.006 0.25 6.65 0.345 ;
      RECT 5.96 0.194 6.006 0.322 ;
      RECT 3.657 0.171 3.797 0.32 ;
      RECT 5.922 0.25 6.65 0.28 ;
      RECT 3.657 0.171 5.96 0.261 ;
      RECT 3.657 0.233 6.039 0.261 ;
      RECT 5.975 0.779 6.115 0.869 ;
      RECT 5.975 0.527 6.065 0.869 ;
      RECT 5.285 0.531 6.065 0.621 ;
      RECT 5.743 0.527 6.065 0.621 ;
      RECT 5.743 0.351 5.883 0.621 ;
      RECT 3.536 1.139 4.862 1.229 ;
      RECT 4.772 0.891 4.862 1.229 ;
      RECT 4.772 0.891 5.245 0.981 ;
      RECT 3.263 1.06 3.403 1.229 ;
      RECT 2.417 1.065 2.557 1.226 ;
      RECT 2.227 1.065 2.63 1.155 ;
      RECT 2.5 1.06 3.403 1.15 ;
      RECT 2.213 1.02 2.227 1.148 ;
      RECT 2.167 0.99 2.213 1.118 ;
      RECT 2.167 1.065 3.434 1.103 ;
      RECT 2.495 1.062 3.472 1.068 ;
      RECT 2.144 1.046 2.265 1.084 ;
      RECT 3.333 1.037 3.472 1.068 ;
      RECT 2.098 0.41 2.167 1.049 ;
      RECT 3.379 1.002 4.37 1.049 ;
      RECT 2.052 0.41 2.167 1.003 ;
      RECT 3.403 0.974 4.412 1.028 ;
      RECT 4.412 0.531 4.458 0.984 ;
      RECT 1.77 0.89 2.167 0.98 ;
      RECT 3.434 0.959 4.458 0.984 ;
      RECT 4.37 0.9 4.412 1.028 ;
      RECT 4.332 0.94 4.458 0.984 ;
      RECT 4.412 0.531 4.502 0.939 ;
      RECT 4.412 0.531 4.909 0.621 ;
      RECT 1.712 0.41 2.167 0.5 ;
      RECT 1.712 0.35 1.852 0.5 ;
      RECT 4.154 0.731 4.294 0.869 ;
      RECT 3.887 0.731 4.322 0.821 ;
      RECT 4.232 0.351 4.322 0.821 ;
      RECT 3.328 0.711 3.944 0.801 ;
      RECT 3.314 0.617 3.328 0.745 ;
      RECT 3.276 0.69 3.415 0.719 ;
      RECT 2.68 0.61 3.314 0.7 ;
      RECT 2.68 0.647 3.374 0.7 ;
      RECT 3.952 0.351 4.322 0.441 ;
      RECT 3.098 0.79 3.238 0.97 ;
      RECT 2.595 0.79 3.238 0.88 ;
      RECT 2.561 0.735 2.595 0.863 ;
      RECT 2.529 0.79 3.238 0.83 ;
      RECT 2.483 0.43 2.561 0.791 ;
      RECT 2.483 0.771 2.633 0.791 ;
      RECT 2.437 0.43 2.561 0.745 ;
      RECT 4.002 0.531 4.142 0.641 ;
      RECT 3.453 0.531 4.142 0.621 ;
      RECT 3.419 0.476 3.453 0.604 ;
      RECT 3.373 0.436 3.419 0.564 ;
      RECT 3.369 0.413 3.373 0.539 ;
      RECT 3.369 0.512 3.491 0.539 ;
      RECT 3.352 0.512 3.491 0.529 ;
      RECT 3.214 0.351 3.369 0.52 ;
      RECT 2.437 0.43 3.373 0.52 ;
      RECT 2.317 0.885 2.457 0.975 ;
      RECT 2.303 0.885 2.457 0.968 ;
      RECT 2.257 0.215 2.347 0.938 ;
      RECT 2.257 0.88 2.402 0.938 ;
      RECT 2.257 0.853 2.393 0.938 ;
      RECT 2.257 0.25 3.076 0.34 ;
      RECT 2.257 0.25 3.155 0.28 ;
      RECT 3.117 0.171 3.567 0.261 ;
      RECT 3.038 0.231 3.567 0.261 ;
      RECT 3.076 0.191 3.117 0.32 ;
      RECT 2.257 0.215 2.411 0.34 ;
      RECT 1.944 1.14 2.084 1.23 ;
      RECT 1.725 1.126 2.059 1.216 ;
      RECT 1.682 1.066 1.725 1.195 ;
      RECT 0.887 1.095 1.28 1.185 ;
      RECT 1.644 1.045 1.682 1.154 ;
      RECT 0.887 1.095 1.33 1.154 ;
      RECT 1.292 1.045 1.682 1.135 ;
      RECT 0.887 1.107 1.763 1.135 ;
      RECT 1.242 1.076 1.725 1.135 ;
      RECT 1.28 1.051 1.292 1.179 ;
      RECT 1.532 0.25 1.622 1.135 ;
      RECT 1.531 0.25 1.622 0.365 ;
      RECT 1.506 0.25 1.622 0.353 ;
      RECT 0.838 0.25 1.622 0.34 ;
      RECT 1.957 0.17 2.097 0.32 ;
      RECT 0.838 0.25 1.674 0.279 ;
      RECT 1.636 0.17 2.097 0.26 ;
      RECT 1.556 0.227 2.097 0.26 ;
      RECT 1.622 0.177 1.636 0.305 ;
      RECT 0.838 0.206 0.978 0.34 ;
      RECT 1.602 0.194 2.097 0.26 ;
      RECT 0.045 1.08 0.271 1.17 ;
      RECT 0.045 0.442 0.135 1.17 ;
      RECT 0.946 0.75 1.261 0.86 ;
      RECT 0.946 0.442 1.036 0.86 ;
      RECT 0.711 0.442 1.036 0.58 ;
      RECT 0.045 0.442 1.036 0.532 ;
      RECT 0.153 0.237 0.243 0.532 ;
  END
END SDFFSRX0P5H7R

MACRO SDFFSRX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRX1H7R 0 0 ;
  SIZE 8.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 8.8 1.48 ;
        RECT 8.065 1.028 8.155 1.48 ;
        RECT 7.35 1.24 7.49 1.48 ;
        RECT 6.386 1.24 6.526 1.48 ;
        RECT 5.385 1.24 5.525 1.48 ;
        RECT 2.807 1.24 2.947 1.48 ;
        RECT 1.466 1.225 1.606 1.48 ;
        RECT 0.381 1.095 0.521 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 8.8 0.08 ;
        RECT 8.065 -0.08 8.155 0.41 ;
        RECT 7.27 -0.08 7.41 0.305 ;
        RECT 6.103 -0.08 6.243 0.16 ;
        RECT 2.86 -0.08 3 0.16 ;
        RECT 1.378 -0.08 1.518 0.16 ;
        RECT 0.378 -0.08 0.518 0.305 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.728 0.59 1.95 0.795 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.622 0.631 0.808 ;
        RECT 0.43 0.622 0.631 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 8.315 0.65 8.575 0.75 ;
        RECT 8.315 0.63 8.563 0.75 ;
        RECT 8.315 0.286 8.405 1.082 ;
      LAYER MET2 ;
        RECT 8.45 0.43 8.55 0.96 ;
      LAYER VIA1 ;
        RECT 8.455 0.655 8.545 0.745 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.705 0.225 7.95 0.375 ;
        RECT 7.705 0.225 7.795 0.945 ;
      LAYER MET2 ;
        RECT 7.85 0.18 7.95 0.56 ;
      LAYER VIA1 ;
        RECT 7.855 0.255 7.945 0.345 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.205 0.45 6.375 0.55 ;
        RECT 6.205 0.45 6.295 0.749 ;
      LAYER MET2 ;
        RECT 6.25 0.225 6.35 0.76 ;
      LAYER VIA1 ;
        RECT 6.255 0.455 6.345 0.545 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.9 0.856 0.99 ;
        RECT 0.766 0.74 0.856 0.99 ;
        RECT 0.225 0.85 0.375 0.99 ;
        RECT 0.225 0.655 0.34 0.99 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.16 0.445 1.442 0.602 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END SI
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.465 0.45 6.775 0.628 ;
      LAYER MET2 ;
        RECT 6.65 0.225 6.75 0.76 ;
      LAYER VIA1 ;
        RECT 6.655 0.455 6.745 0.545 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 5.615 1.14 6.267 1.23 ;
      RECT 4.952 1.071 5.092 1.229 ;
      RECT 5.615 1.14 6.308 1.21 ;
      RECT 5.615 1.14 6.347 1.17 ;
      RECT 4.952 1.071 5.34 1.161 ;
      RECT 7.885 0.546 7.975 1.15 ;
      RECT 5.295 1.059 5.705 1.149 ;
      RECT 6.228 1.12 7.975 1.15 ;
      RECT 7.525 1.059 7.975 1.15 ;
      RECT 6.267 1.08 7.975 1.15 ;
      RECT 6.308 1.06 7.975 1.15 ;
      RECT 7.525 0.395 7.615 1.15 ;
      RECT 7.885 0.546 8.176 0.636 ;
      RECT 7.02 0.395 7.615 0.485 ;
      RECT 7.02 0.264 7.16 0.485 ;
      RECT 5.795 0.959 6.191 1.049 ;
      RECT 5.795 0.959 6.232 1.029 ;
      RECT 4.592 0.711 4.682 0.997 ;
      RECT 5.795 0.959 6.27 0.989 ;
      RECT 6.865 0.575 6.955 0.97 ;
      RECT 6.153 0.94 6.955 0.97 ;
      RECT 6.232 0.88 6.955 0.97 ;
      RECT 5.795 0.711 5.885 1.049 ;
      RECT 6.191 0.9 6.955 0.97 ;
      RECT 4.592 0.711 5.885 0.801 ;
      RECT 6.865 0.575 7.247 0.715 ;
      RECT 4.999 0.351 5.089 0.801 ;
      RECT 4.513 0.351 5.623 0.441 ;
      RECT 6.001 0.25 6.65 0.34 ;
      RECT 5.96 0.191 6.001 0.32 ;
      RECT 3.657 0.171 3.797 0.32 ;
      RECT 5.922 0.25 6.65 0.28 ;
      RECT 3.657 0.171 5.96 0.261 ;
      RECT 3.657 0.231 6.039 0.261 ;
      RECT 5.975 0.779 6.115 0.869 ;
      RECT 5.975 0.527 6.065 0.869 ;
      RECT 5.285 0.531 6.065 0.621 ;
      RECT 5.743 0.527 6.065 0.621 ;
      RECT 5.743 0.351 5.883 0.621 ;
      RECT 3.536 1.139 4.862 1.229 ;
      RECT 4.772 0.891 4.862 1.229 ;
      RECT 4.772 0.891 5.245 0.981 ;
      RECT 3.263 1.06 3.403 1.229 ;
      RECT 2.417 1.065 2.557 1.226 ;
      RECT 2.227 1.065 2.63 1.155 ;
      RECT 2.5 1.06 3.403 1.15 ;
      RECT 2.213 1.02 2.227 1.148 ;
      RECT 2.167 0.99 2.213 1.118 ;
      RECT 2.167 1.065 3.434 1.103 ;
      RECT 2.495 1.062 3.472 1.068 ;
      RECT 2.144 1.046 2.265 1.084 ;
      RECT 3.333 1.037 3.472 1.068 ;
      RECT 2.098 0.41 2.167 1.049 ;
      RECT 3.379 1.002 4.37 1.049 ;
      RECT 2.052 0.41 2.167 1.003 ;
      RECT 3.403 0.974 4.412 1.028 ;
      RECT 4.412 0.531 4.458 0.984 ;
      RECT 1.77 0.89 2.167 0.98 ;
      RECT 3.434 0.959 4.458 0.984 ;
      RECT 4.37 0.9 4.412 1.028 ;
      RECT 4.332 0.94 4.458 0.984 ;
      RECT 4.412 0.531 4.502 0.939 ;
      RECT 4.412 0.531 4.909 0.621 ;
      RECT 1.712 0.41 2.167 0.5 ;
      RECT 1.712 0.35 1.852 0.5 ;
      RECT 4.154 0.731 4.294 0.869 ;
      RECT 3.887 0.731 4.322 0.821 ;
      RECT 4.232 0.351 4.322 0.821 ;
      RECT 3.328 0.711 3.944 0.801 ;
      RECT 3.314 0.617 3.328 0.745 ;
      RECT 3.276 0.69 3.415 0.719 ;
      RECT 2.68 0.61 3.314 0.7 ;
      RECT 2.68 0.647 3.374 0.7 ;
      RECT 3.952 0.351 4.322 0.441 ;
      RECT 3.098 0.79 3.238 0.97 ;
      RECT 2.595 0.79 3.238 0.88 ;
      RECT 2.561 0.735 2.595 0.863 ;
      RECT 2.529 0.79 3.238 0.83 ;
      RECT 2.483 0.43 2.561 0.791 ;
      RECT 2.483 0.771 2.633 0.791 ;
      RECT 2.437 0.43 2.561 0.745 ;
      RECT 4.002 0.531 4.142 0.641 ;
      RECT 3.453 0.531 4.142 0.621 ;
      RECT 3.419 0.476 3.453 0.604 ;
      RECT 3.373 0.436 3.419 0.564 ;
      RECT 3.369 0.413 3.373 0.539 ;
      RECT 3.369 0.512 3.491 0.539 ;
      RECT 3.352 0.512 3.491 0.529 ;
      RECT 3.214 0.351 3.369 0.52 ;
      RECT 2.437 0.43 3.373 0.52 ;
      RECT 2.317 0.885 2.457 0.975 ;
      RECT 2.303 0.885 2.457 0.968 ;
      RECT 2.257 0.215 2.347 0.938 ;
      RECT 2.257 0.88 2.402 0.938 ;
      RECT 2.257 0.853 2.393 0.938 ;
      RECT 2.257 0.25 3.076 0.34 ;
      RECT 2.257 0.25 3.155 0.28 ;
      RECT 3.117 0.171 3.567 0.261 ;
      RECT 3.038 0.231 3.567 0.261 ;
      RECT 3.076 0.191 3.117 0.32 ;
      RECT 2.257 0.215 2.411 0.34 ;
      RECT 1.739 1.14 2.084 1.23 ;
      RECT 1.728 1.096 1.739 1.225 ;
      RECT 1.682 1.068 1.728 1.196 ;
      RECT 0.887 1.095 1.28 1.185 ;
      RECT 0.887 1.095 1.33 1.154 ;
      RECT 1.644 1.126 2.059 1.154 ;
      RECT 1.292 1.045 1.682 1.135 ;
      RECT 0.887 1.114 1.763 1.135 ;
      RECT 1.242 1.076 1.728 1.135 ;
      RECT 1.28 1.051 1.292 1.179 ;
      RECT 1.532 0.25 1.622 1.135 ;
      RECT 1.531 0.25 1.622 0.365 ;
      RECT 1.506 0.25 1.622 0.353 ;
      RECT 0.838 0.25 1.622 0.34 ;
      RECT 1.957 0.17 2.097 0.32 ;
      RECT 0.838 0.25 1.674 0.279 ;
      RECT 1.636 0.17 2.097 0.26 ;
      RECT 1.556 0.227 2.097 0.26 ;
      RECT 1.622 0.177 1.636 0.305 ;
      RECT 0.838 0.206 0.978 0.34 ;
      RECT 1.602 0.194 2.097 0.26 ;
      RECT 0.045 1.08 0.271 1.17 ;
      RECT 0.045 0.442 0.135 1.17 ;
      RECT 0.946 0.75 1.261 0.86 ;
      RECT 0.946 0.442 1.036 0.86 ;
      RECT 0.711 0.442 1.036 0.58 ;
      RECT 0.045 0.442 1.036 0.532 ;
      RECT 0.153 0.237 0.243 0.532 ;
  END
END SDFFSRX1H7R

MACRO SDFFSRX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRX2H7R 0 0 ;
  SIZE 8.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 8.8 1.48 ;
        RECT 8.065 1.028 8.155 1.48 ;
        RECT 7.35 1.24 7.49 1.48 ;
        RECT 6.386 1.24 6.526 1.48 ;
        RECT 5.385 1.24 5.525 1.48 ;
        RECT 2.807 1.24 2.947 1.48 ;
        RECT 1.466 1.225 1.606 1.48 ;
        RECT 0.381 1.095 0.521 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 8.8 0.08 ;
        RECT 8.065 -0.08 8.155 0.33 ;
        RECT 7.27 -0.08 7.41 0.305 ;
        RECT 6.103 -0.08 6.243 0.16 ;
        RECT 2.86 -0.08 3 0.16 ;
        RECT 1.378 -0.08 1.518 0.16 ;
        RECT 0.378 -0.08 0.518 0.305 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 1.728 0.59 1.95 0.795 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.455 0.622 0.631 0.808 ;
        RECT 0.43 0.622 0.631 0.775 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 8.315 0.63 8.575 0.75 ;
        RECT 8.315 0.286 8.405 1.082 ;
      LAYER MET2 ;
        RECT 8.45 0.43 8.55 0.96 ;
      LAYER VIA1 ;
        RECT 8.455 0.655 8.545 0.745 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.705 0.225 7.95 0.375 ;
        RECT 7.705 0.225 7.795 0.945 ;
      LAYER MET2 ;
        RECT 7.85 0.18 7.95 0.56 ;
      LAYER VIA1 ;
        RECT 7.855 0.255 7.945 0.345 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.205 0.45 6.375 0.55 ;
        RECT 6.205 0.45 6.295 0.749 ;
      LAYER MET2 ;
        RECT 6.25 0.225 6.35 0.76 ;
      LAYER VIA1 ;
        RECT 6.255 0.455 6.345 0.545 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.9 0.856 0.99 ;
        RECT 0.766 0.74 0.856 0.99 ;
        RECT 0.225 0.85 0.375 0.99 ;
        RECT 0.225 0.655 0.34 0.99 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.16 0.445 1.442 0.602 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END SI
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.465 0.455 6.775 0.628 ;
        RECT 6.625 0.45 6.775 0.628 ;
      LAYER MET2 ;
        RECT 6.65 0.225 6.75 0.76 ;
      LAYER VIA1 ;
        RECT 6.655 0.455 6.745 0.545 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 5.615 1.14 6.267 1.23 ;
      RECT 4.952 1.071 5.092 1.229 ;
      RECT 5.615 1.14 6.308 1.21 ;
      RECT 5.615 1.14 6.347 1.17 ;
      RECT 4.952 1.071 5.335 1.161 ;
      RECT 7.885 0.546 7.975 1.15 ;
      RECT 5.29 1.059 5.705 1.149 ;
      RECT 6.228 1.12 7.975 1.15 ;
      RECT 7.525 1.059 7.975 1.15 ;
      RECT 6.267 1.08 7.975 1.15 ;
      RECT 6.308 1.06 7.975 1.15 ;
      RECT 7.525 0.395 7.615 1.15 ;
      RECT 7.885 0.546 8.176 0.636 ;
      RECT 7.02 0.395 7.615 0.485 ;
      RECT 7.02 0.264 7.16 0.485 ;
      RECT 5.795 0.959 6.191 1.049 ;
      RECT 5.795 0.959 6.232 1.029 ;
      RECT 4.592 0.711 4.682 0.997 ;
      RECT 5.795 0.959 6.27 0.989 ;
      RECT 6.865 0.575 6.955 0.97 ;
      RECT 6.153 0.94 6.955 0.97 ;
      RECT 6.232 0.88 6.955 0.97 ;
      RECT 5.795 0.711 5.885 1.049 ;
      RECT 6.191 0.9 6.955 0.97 ;
      RECT 4.592 0.711 5.885 0.801 ;
      RECT 6.865 0.575 7.247 0.715 ;
      RECT 4.999 0.351 5.089 0.801 ;
      RECT 4.513 0.351 5.623 0.441 ;
      RECT 6.001 0.25 6.65 0.34 ;
      RECT 5.96 0.191 6.001 0.32 ;
      RECT 3.657 0.171 3.797 0.32 ;
      RECT 5.922 0.25 6.65 0.28 ;
      RECT 3.657 0.171 5.96 0.261 ;
      RECT 3.657 0.231 6.039 0.261 ;
      RECT 5.975 0.779 6.115 0.869 ;
      RECT 5.975 0.527 6.065 0.869 ;
      RECT 5.285 0.531 6.065 0.621 ;
      RECT 5.743 0.527 6.065 0.621 ;
      RECT 5.743 0.351 5.883 0.621 ;
      RECT 3.536 1.139 4.862 1.229 ;
      RECT 4.772 0.891 4.862 1.229 ;
      RECT 4.772 0.891 5.245 0.981 ;
      RECT 3.263 1.06 3.403 1.229 ;
      RECT 2.417 1.065 2.557 1.226 ;
      RECT 2.227 1.065 2.63 1.155 ;
      RECT 2.5 1.06 3.403 1.15 ;
      RECT 2.213 1.02 2.227 1.148 ;
      RECT 2.167 0.99 2.213 1.118 ;
      RECT 2.167 1.065 3.434 1.103 ;
      RECT 2.495 1.062 3.472 1.068 ;
      RECT 2.144 1.046 2.265 1.084 ;
      RECT 3.333 1.037 3.472 1.068 ;
      RECT 2.098 0.41 2.167 1.049 ;
      RECT 3.379 1.002 4.37 1.049 ;
      RECT 2.052 0.41 2.167 1.003 ;
      RECT 3.403 0.974 4.412 1.028 ;
      RECT 4.412 0.531 4.458 0.984 ;
      RECT 1.77 0.89 2.167 0.98 ;
      RECT 3.434 0.959 4.458 0.984 ;
      RECT 4.37 0.9 4.412 1.028 ;
      RECT 4.332 0.94 4.458 0.984 ;
      RECT 4.412 0.531 4.502 0.939 ;
      RECT 4.412 0.531 4.909 0.621 ;
      RECT 1.712 0.41 2.167 0.5 ;
      RECT 1.712 0.35 1.852 0.5 ;
      RECT 4.154 0.731 4.294 0.869 ;
      RECT 3.887 0.731 4.322 0.821 ;
      RECT 4.232 0.351 4.322 0.821 ;
      RECT 3.328 0.711 3.944 0.801 ;
      RECT 3.314 0.617 3.328 0.745 ;
      RECT 3.276 0.69 3.415 0.719 ;
      RECT 2.68 0.61 3.314 0.7 ;
      RECT 2.68 0.647 3.374 0.7 ;
      RECT 3.952 0.351 4.322 0.441 ;
      RECT 3.098 0.79 3.238 0.97 ;
      RECT 2.595 0.79 3.238 0.88 ;
      RECT 2.561 0.735 2.595 0.863 ;
      RECT 2.517 0.771 2.633 0.824 ;
      RECT 2.471 0.43 2.561 0.779 ;
      RECT 4.002 0.531 4.142 0.641 ;
      RECT 2.437 0.43 2.561 0.624 ;
      RECT 3.453 0.531 4.142 0.621 ;
      RECT 3.419 0.476 3.453 0.604 ;
      RECT 3.373 0.436 3.419 0.564 ;
      RECT 3.369 0.413 3.373 0.539 ;
      RECT 3.369 0.512 3.491 0.539 ;
      RECT 3.352 0.512 3.491 0.529 ;
      RECT 3.214 0.351 3.369 0.52 ;
      RECT 2.437 0.43 3.373 0.52 ;
      RECT 2.317 0.885 2.457 0.975 ;
      RECT 2.303 0.885 2.457 0.968 ;
      RECT 2.257 0.215 2.347 0.938 ;
      RECT 2.257 0.88 2.402 0.938 ;
      RECT 2.257 0.853 2.393 0.938 ;
      RECT 2.257 0.25 3.076 0.34 ;
      RECT 2.257 0.25 3.155 0.28 ;
      RECT 3.117 0.171 3.567 0.261 ;
      RECT 3.038 0.231 3.567 0.261 ;
      RECT 3.076 0.191 3.117 0.32 ;
      RECT 2.257 0.215 2.411 0.34 ;
      RECT 1.944 1.14 2.084 1.23 ;
      RECT 1.725 1.126 2.059 1.216 ;
      RECT 1.682 1.066 1.725 1.195 ;
      RECT 0.887 1.095 1.28 1.185 ;
      RECT 1.644 1.045 1.682 1.154 ;
      RECT 0.887 1.095 1.33 1.154 ;
      RECT 1.292 1.045 1.682 1.135 ;
      RECT 0.887 1.107 1.763 1.135 ;
      RECT 1.242 1.076 1.725 1.135 ;
      RECT 1.28 1.051 1.292 1.179 ;
      RECT 1.532 0.25 1.622 1.135 ;
      RECT 1.531 0.25 1.622 0.365 ;
      RECT 1.506 0.25 1.622 0.353 ;
      RECT 0.838 0.25 1.622 0.34 ;
      RECT 1.957 0.17 2.097 0.32 ;
      RECT 0.838 0.25 1.674 0.279 ;
      RECT 1.636 0.17 2.097 0.26 ;
      RECT 1.556 0.227 2.097 0.26 ;
      RECT 1.622 0.177 1.636 0.305 ;
      RECT 0.838 0.206 0.978 0.34 ;
      RECT 1.602 0.194 2.097 0.26 ;
      RECT 0.045 1.08 0.271 1.17 ;
      RECT 0.045 0.442 0.135 1.17 ;
      RECT 0.946 0.75 1.261 0.86 ;
      RECT 0.946 0.442 1.036 0.86 ;
      RECT 0.711 0.442 1.036 0.58 ;
      RECT 0.045 0.442 1.036 0.532 ;
      RECT 0.153 0.237 0.243 0.532 ;
  END
END SDFFSRX2H7R

MACRO SDFFSX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSX0P5H7R 0 0 ;
  SIZE 8.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 8.2 1.48 ;
        RECT 7.57 1.07 7.66 1.48 ;
        RECT 6.85 1.07 6.94 1.48 ;
        RECT 5.83 0.98 5.92 1.48 ;
        RECT 3.745 1.125 3.885 1.48 ;
        RECT 3.045 1.24 3.185 1.48 ;
        RECT 1.595 1.07 1.685 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 8.2 0.08 ;
        RECT 7.26 -0.08 7.35 0.35 ;
        RECT 6.645 -0.08 6.735 0.35 ;
        RECT 6.165 -0.08 6.255 0.35 ;
        RECT 3.04 -0.08 3.18 0.16 ;
        RECT 1.595 -0.08 1.685 0.35 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 4.155 0.835 4.405 1.04 ;
      LAYER MET2 ;
        RECT 4.25 0.625 4.35 1.16 ;
      LAYER VIA1 ;
        RECT 4.255 0.855 4.345 0.945 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.56 0.595 0.65 ;
        RECT 0.225 0.45 0.375 0.65 ;
      LAYER MET2 ;
        RECT 0.25 0.18 0.35 0.585 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.82 1.055 7.945 1.195 ;
        RECT 7.845 0.395 7.945 1.195 ;
        RECT 7.51 0.395 7.945 0.485 ;
        RECT 7.51 0.21 7.6 0.485 ;
      LAYER MET2 ;
        RECT 7.85 0.84 7.95 1.22 ;
      LAYER VIA1 ;
        RECT 7.855 1.055 7.945 1.145 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.21 0.655 7.3 1.05 ;
        RECT 7.03 0.655 7.3 0.745 ;
        RECT 7.03 0.21 7.145 0.745 ;
      LAYER MET2 ;
        RECT 7.05 0.18 7.15 0.56 ;
      LAYER VIA1 ;
        RECT 7.055 0.255 7.145 0.345 ;
    END
  END QN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.74 0.855 0.855 ;
        RECT 0.225 0.74 0.375 0.95 ;
      LAYER MET2 ;
        RECT 0.25 0.815 0.35 1.22 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.595 0.455 1.788 0.61 ;
      LAYER MET2 ;
        RECT 1.65 0.23 1.75 0.76 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END SI
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.255 0.62 6.4 0.82 ;
      LAYER MET2 ;
        RECT 6.25 0.425 6.35 0.96 ;
      LAYER VIA1 ;
        RECT 6.255 0.655 6.345 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 7.03 1.14 7.48 1.23 ;
      RECT 7.39 0.575 7.48 1.23 ;
      RECT 7.03 0.89 7.12 1.23 ;
      RECT 6.37 0.91 6.58 1 ;
      RECT 6.49 0.44 6.58 1 ;
      RECT 6.85 0.89 7.12 0.98 ;
      RECT 6.85 0.44 6.94 0.98 ;
      RECT 5.835 0.53 5.925 0.71 ;
      RECT 7.39 0.575 7.755 0.665 ;
      RECT 5.835 0.53 6.155 0.62 ;
      RECT 6.065 0.44 6.94 0.53 ;
      RECT 6.395 0.255 6.485 0.53 ;
      RECT 6.19 1.14 6.76 1.23 ;
      RECT 6.67 0.68 6.76 1.23 ;
      RECT 6.19 0.99 6.28 1.23 ;
      RECT 6.01 0.99 6.28 1.08 ;
      RECT 5.12 0.35 5.21 0.995 ;
      RECT 6.01 0.8 6.1 1.08 ;
      RECT 5.655 0.8 6.1 0.89 ;
      RECT 5.655 0.35 5.745 0.89 ;
      RECT 4.715 0.35 5.745 0.44 ;
      RECT 3.64 0.35 4.365 0.44 ;
      RECT 4.275 0.17 4.365 0.44 ;
      RECT 5.835 0.325 5.975 0.415 ;
      RECT 5.835 0.17 5.925 0.415 ;
      RECT 4.275 0.17 5.925 0.26 ;
      RECT 3.975 1.14 5.415 1.23 ;
      RECT 5.325 0.61 5.415 1.23 ;
      RECT 3.975 0.945 4.065 1.23 ;
      RECT 3.4 0.88 3.49 1.05 ;
      RECT 3.4 0.945 4.065 1.035 ;
      RECT 2.63 0.88 3.49 0.97 ;
      RECT 2.63 0.498 2.72 0.97 ;
      RECT 5.325 0.61 5.565 0.7 ;
      RECT 2.63 0.498 2.721 0.559 ;
      RECT 2.63 0.498 2.759 0.539 ;
      RECT 2.63 0.498 3.334 0.52 ;
      RECT 2.676 0.453 3.376 0.499 ;
      RECT 2.72 0.43 3.414 0.459 ;
      RECT 3.334 0.371 3.376 0.499 ;
      RECT 3.376 0.35 3.52 0.44 ;
      RECT 3.296 0.411 3.52 0.44 ;
      RECT 4.505 0.93 4.875 1.02 ;
      RECT 4.505 0.35 4.595 1.02 ;
      RECT 2.865 0.61 4.595 0.7 ;
      RECT 4.455 0.35 4.595 0.44 ;
      RECT 1.955 0.17 2.045 1.05 ;
      RECT 1.955 0.66 2.125 0.8 ;
      RECT 2.86 0.25 3.258 0.34 ;
      RECT 2.86 0.25 3.338 0.279 ;
      RECT 3.3 0.17 4.185 0.26 ;
      RECT 3.22 0.231 4.185 0.26 ;
      RECT 3.258 0.191 3.3 0.319 ;
      RECT 1.955 0.17 2.95 0.26 ;
      RECT 3.305 1.14 3.655 1.23 ;
      RECT 2.45 1.14 2.927 1.23 ;
      RECT 3.263 1.14 3.655 1.209 ;
      RECT 2.45 1.14 2.969 1.209 ;
      RECT 3.225 1.14 3.655 1.169 ;
      RECT 2.45 1.14 3.007 1.169 ;
      RECT 2.969 1.06 3.263 1.15 ;
      RECT 2.889 1.121 3.343 1.15 ;
      RECT 2.45 0.35 2.54 1.23 ;
      RECT 2.927 1.081 3.305 1.15 ;
      RECT 2.425 0.35 2.565 0.44 ;
      RECT 1.775 1.14 2.29 1.23 ;
      RECT 0.785 1.05 1.505 1.14 ;
      RECT 1.415 0.25 1.505 1.14 ;
      RECT 2.2 0.89 2.29 1.23 ;
      RECT 1.775 0.89 1.865 1.23 ;
      RECT 2.215 0.35 2.305 0.98 ;
      RECT 1.415 0.89 1.865 0.98 ;
      RECT 2.175 0.35 2.315 0.44 ;
      RECT 0.865 0.25 1.505 0.34 ;
      RECT 0.045 1.05 0.185 1.14 ;
      RECT 0.045 0.25 0.135 1.14 ;
      RECT 0.945 0.795 1.325 0.885 ;
      RECT 0.945 0.495 1.035 0.885 ;
      RECT 0.685 0.495 1.035 0.585 ;
      RECT 0.685 0.265 0.775 0.585 ;
      RECT 0.045 0.265 0.775 0.355 ;
      RECT 0.045 0.25 0.185 0.355 ;
  END
END SDFFSX0P5H7R

MACRO SDFFSX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSX1H7R 0 0 ;
  SIZE 8.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 8.2 1.48 ;
        RECT 7.57 1.07 7.66 1.48 ;
        RECT 6.85 1.07 6.94 1.48 ;
        RECT 5.83 0.98 5.92 1.48 ;
        RECT 3.745 1.125 3.885 1.48 ;
        RECT 3.045 1.24 3.185 1.48 ;
        RECT 1.595 1.07 1.685 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 8.2 0.08 ;
        RECT 7.26 -0.08 7.35 0.35 ;
        RECT 6.645 -0.08 6.735 0.35 ;
        RECT 6.165 -0.08 6.255 0.35 ;
        RECT 3.04 -0.08 3.18 0.16 ;
        RECT 1.595 -0.08 1.685 0.35 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 4.155 0.835 4.405 1.04 ;
      LAYER MET2 ;
        RECT 4.25 0.625 4.35 1.16 ;
      LAYER VIA1 ;
        RECT 4.255 0.855 4.345 0.945 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.56 0.595 0.65 ;
        RECT 0.225 0.45 0.376 0.65 ;
      LAYER MET2 ;
        RECT 0.25 0.18 0.35 0.585 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.82 1.02 7.945 1.195 ;
        RECT 7.845 0.395 7.935 1.195 ;
        RECT 7.51 0.395 7.935 0.485 ;
        RECT 7.51 0.21 7.6 0.485 ;
      LAYER MET2 ;
        RECT 7.85 0.84 7.95 1.22 ;
      LAYER VIA1 ;
        RECT 7.855 1.055 7.945 1.145 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.21 0.655 7.3 1.05 ;
        RECT 7.03 0.655 7.3 0.745 ;
        RECT 7.03 0.21 7.145 0.745 ;
      LAYER MET2 ;
        RECT 7.05 0.18 7.15 0.56 ;
      LAYER VIA1 ;
        RECT 7.055 0.255 7.145 0.345 ;
    END
  END QN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.74 0.855 0.855 ;
        RECT 0.225 0.74 0.375 0.95 ;
      LAYER MET2 ;
        RECT 0.25 0.815 0.35 1.22 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.595 0.455 1.788 0.61 ;
      LAYER MET2 ;
        RECT 1.65 0.23 1.75 0.76 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END SI
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.255 0.62 6.4 0.82 ;
      LAYER MET2 ;
        RECT 6.25 0.425 6.35 0.96 ;
      LAYER VIA1 ;
        RECT 6.255 0.655 6.345 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 7.03 1.14 7.48 1.23 ;
      RECT 7.39 0.575 7.48 1.23 ;
      RECT 7.03 0.89 7.12 1.23 ;
      RECT 6.37 0.91 6.58 1 ;
      RECT 6.49 0.44 6.58 1 ;
      RECT 6.85 0.89 7.12 0.98 ;
      RECT 6.85 0.44 6.94 0.98 ;
      RECT 5.835 0.53 5.925 0.71 ;
      RECT 7.39 0.575 7.755 0.665 ;
      RECT 5.835 0.53 6.155 0.62 ;
      RECT 6.065 0.44 6.94 0.53 ;
      RECT 6.395 0.275 6.485 0.53 ;
      RECT 6.19 1.14 6.76 1.23 ;
      RECT 6.67 0.68 6.76 1.23 ;
      RECT 6.19 0.99 6.28 1.23 ;
      RECT 6.01 0.99 6.28 1.08 ;
      RECT 5.12 0.35 5.21 0.995 ;
      RECT 6.01 0.8 6.1 1.08 ;
      RECT 5.655 0.8 6.1 0.89 ;
      RECT 5.655 0.35 5.745 0.89 ;
      RECT 4.715 0.35 5.745 0.44 ;
      RECT 5.835 0.35 5.975 0.44 ;
      RECT 3.64 0.35 4.365 0.44 ;
      RECT 4.275 0.17 4.365 0.44 ;
      RECT 5.835 0.17 5.925 0.44 ;
      RECT 4.275 0.17 5.925 0.26 ;
      RECT 3.975 1.14 5.415 1.23 ;
      RECT 5.325 0.61 5.415 1.23 ;
      RECT 3.975 0.945 4.065 1.23 ;
      RECT 3.4 0.88 3.49 1.05 ;
      RECT 3.4 0.945 4.065 1.035 ;
      RECT 2.63 0.88 3.49 0.97 ;
      RECT 2.63 0.498 2.72 0.97 ;
      RECT 5.325 0.61 5.565 0.7 ;
      RECT 2.63 0.498 2.721 0.559 ;
      RECT 2.63 0.498 2.759 0.539 ;
      RECT 2.63 0.498 3.334 0.52 ;
      RECT 2.676 0.453 3.376 0.499 ;
      RECT 2.72 0.43 3.414 0.459 ;
      RECT 3.334 0.371 3.376 0.499 ;
      RECT 3.376 0.35 3.52 0.44 ;
      RECT 3.296 0.411 3.52 0.44 ;
      RECT 4.505 0.91 4.875 1 ;
      RECT 4.505 0.35 4.595 1 ;
      RECT 2.865 0.61 4.595 0.7 ;
      RECT 4.455 0.35 4.595 0.44 ;
      RECT 1.955 0.17 2.045 1.05 ;
      RECT 1.955 0.66 2.125 0.8 ;
      RECT 2.86 0.25 3.258 0.34 ;
      RECT 2.86 0.25 3.338 0.279 ;
      RECT 3.3 0.17 4.185 0.26 ;
      RECT 3.22 0.231 4.185 0.26 ;
      RECT 3.258 0.191 3.3 0.319 ;
      RECT 1.955 0.17 2.95 0.26 ;
      RECT 3.305 1.14 3.655 1.23 ;
      RECT 2.45 1.14 2.927 1.23 ;
      RECT 3.263 1.14 3.655 1.209 ;
      RECT 2.45 1.14 2.969 1.209 ;
      RECT 3.225 1.14 3.655 1.169 ;
      RECT 2.45 1.14 3.007 1.169 ;
      RECT 2.969 1.06 3.263 1.15 ;
      RECT 2.889 1.121 3.343 1.15 ;
      RECT 2.45 0.35 2.54 1.23 ;
      RECT 2.927 1.081 3.305 1.15 ;
      RECT 2.425 0.35 2.565 0.44 ;
      RECT 1.775 1.14 2.315 1.23 ;
      RECT 2.215 0.35 2.315 1.23 ;
      RECT 0.785 1.05 1.505 1.14 ;
      RECT 1.415 0.25 1.505 1.14 ;
      RECT 2.2 0.89 2.315 1.23 ;
      RECT 1.775 0.89 1.865 1.23 ;
      RECT 1.415 0.89 1.865 0.98 ;
      RECT 2.175 0.35 2.315 0.44 ;
      RECT 0.865 0.25 1.505 0.34 ;
      RECT 0.045 1.05 0.185 1.14 ;
      RECT 0.045 0.25 0.135 1.14 ;
      RECT 0.945 0.795 1.325 0.885 ;
      RECT 0.945 0.495 1.035 0.885 ;
      RECT 0.685 0.495 1.035 0.585 ;
      RECT 0.685 0.265 0.775 0.585 ;
      RECT 0.045 0.265 0.775 0.355 ;
      RECT 0.045 0.25 0.185 0.355 ;
  END
END SDFFSX1H7R

MACRO SDFFSX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSX2H7R 0 0 ;
  SIZE 8.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 8.2 1.48 ;
        RECT 7.57 1.07 7.66 1.48 ;
        RECT 6.85 1.07 6.94 1.48 ;
        RECT 5.83 0.98 5.92 1.48 ;
        RECT 3.745 1.125 3.885 1.48 ;
        RECT 3.045 1.24 3.185 1.48 ;
        RECT 1.595 1.07 1.685 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 8.2 0.08 ;
        RECT 7.26 -0.08 7.35 0.35 ;
        RECT 6.645 -0.08 6.735 0.35 ;
        RECT 6.165 -0.08 6.255 0.35 ;
        RECT 3.04 -0.08 3.18 0.16 ;
        RECT 1.595 -0.08 1.685 0.35 ;
        RECT 0.31 -0.08 0.45 0.175 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 4.155 0.835 4.405 1.04 ;
      LAYER MET2 ;
        RECT 4.25 0.625 4.35 1.16 ;
      LAYER VIA1 ;
        RECT 4.255 0.855 4.345 0.945 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.56 0.595 0.65 ;
        RECT 0.225 0.45 0.375 0.65 ;
      LAYER MET2 ;
        RECT 0.25 0.18 0.35 0.585 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.82 0.855 7.945 1.195 ;
        RECT 7.845 0.395 7.945 1.195 ;
        RECT 7.51 0.395 7.945 0.485 ;
        RECT 7.51 0.21 7.6 0.485 ;
      LAYER MET2 ;
        RECT 7.85 0.84 7.95 1.22 ;
      LAYER VIA1 ;
        RECT 7.855 1.055 7.945 1.145 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.21 0.655 7.3 1.05 ;
        RECT 7.03 0.655 7.3 0.745 ;
        RECT 7.03 0.21 7.145 0.745 ;
      LAYER MET2 ;
        RECT 7.05 0.18 7.15 0.56 ;
      LAYER VIA1 ;
        RECT 7.055 0.255 7.145 0.345 ;
    END
  END QN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.74 0.855 0.855 ;
        RECT 0.225 0.74 0.375 0.95 ;
      LAYER MET2 ;
        RECT 0.25 0.815 0.35 1.22 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.595 0.455 1.788 0.61 ;
      LAYER MET2 ;
        RECT 1.65 0.23 1.75 0.76 ;
      LAYER VIA1 ;
        RECT 1.655 0.455 1.745 0.545 ;
    END
  END SI
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.255 0.62 6.4 0.82 ;
      LAYER MET2 ;
        RECT 6.25 0.425 6.35 0.96 ;
      LAYER VIA1 ;
        RECT 6.255 0.655 6.345 0.745 ;
    END
  END SN
  OBS
    LAYER MET1 ;
      RECT 7.03 1.14 7.48 1.23 ;
      RECT 7.39 0.575 7.48 1.23 ;
      RECT 7.03 0.89 7.12 1.23 ;
      RECT 6.37 0.91 6.58 1 ;
      RECT 6.49 0.44 6.58 1 ;
      RECT 6.85 0.89 7.12 0.98 ;
      RECT 6.85 0.44 6.94 0.98 ;
      RECT 5.835 0.53 5.925 0.71 ;
      RECT 7.39 0.575 7.755 0.665 ;
      RECT 5.835 0.53 6.155 0.62 ;
      RECT 6.065 0.44 6.94 0.53 ;
      RECT 6.395 0.295 6.485 0.53 ;
      RECT 6.19 1.14 6.76 1.23 ;
      RECT 6.67 0.68 6.76 1.23 ;
      RECT 6.19 0.99 6.28 1.23 ;
      RECT 6.01 0.99 6.28 1.08 ;
      RECT 5.12 0.35 5.21 0.995 ;
      RECT 6.01 0.8 6.1 1.08 ;
      RECT 5.655 0.8 6.1 0.89 ;
      RECT 5.655 0.35 5.745 0.89 ;
      RECT 4.715 0.35 5.745 0.44 ;
      RECT 5.835 0.35 5.975 0.44 ;
      RECT 3.64 0.35 4.365 0.44 ;
      RECT 4.275 0.17 4.365 0.44 ;
      RECT 5.835 0.17 5.925 0.44 ;
      RECT 4.275 0.17 5.925 0.26 ;
      RECT 3.975 1.14 5.415 1.23 ;
      RECT 5.325 0.61 5.415 1.23 ;
      RECT 3.975 0.945 4.065 1.23 ;
      RECT 3.4 0.88 3.49 1.05 ;
      RECT 3.4 0.945 4.065 1.035 ;
      RECT 2.63 0.88 3.49 0.97 ;
      RECT 2.63 0.498 2.72 0.97 ;
      RECT 5.325 0.61 5.565 0.7 ;
      RECT 2.63 0.498 2.721 0.559 ;
      RECT 2.63 0.498 2.759 0.539 ;
      RECT 2.63 0.498 3.334 0.52 ;
      RECT 2.676 0.453 3.376 0.499 ;
      RECT 2.72 0.43 3.414 0.459 ;
      RECT 3.334 0.371 3.376 0.499 ;
      RECT 3.376 0.35 3.52 0.44 ;
      RECT 3.296 0.411 3.52 0.44 ;
      RECT 4.505 0.88 4.875 0.97 ;
      RECT 4.505 0.35 4.595 0.97 ;
      RECT 2.865 0.61 4.595 0.7 ;
      RECT 4.455 0.35 4.595 0.7 ;
      RECT 1.955 0.17 2.045 1.05 ;
      RECT 1.955 0.66 2.125 0.8 ;
      RECT 2.86 0.25 3.258 0.34 ;
      RECT 2.86 0.25 3.338 0.279 ;
      RECT 3.3 0.17 4.185 0.26 ;
      RECT 3.22 0.231 4.185 0.26 ;
      RECT 3.258 0.191 3.3 0.319 ;
      RECT 1.955 0.17 2.95 0.26 ;
      RECT 3.305 1.14 3.655 1.23 ;
      RECT 2.45 1.14 2.927 1.23 ;
      RECT 3.263 1.14 3.655 1.209 ;
      RECT 2.45 1.14 2.969 1.209 ;
      RECT 3.225 1.14 3.655 1.169 ;
      RECT 2.45 1.14 3.007 1.169 ;
      RECT 2.969 1.06 3.263 1.15 ;
      RECT 2.889 1.121 3.343 1.15 ;
      RECT 2.45 0.35 2.54 1.23 ;
      RECT 2.927 1.081 3.305 1.15 ;
      RECT 2.425 0.35 2.565 0.44 ;
      RECT 1.775 1.14 2.315 1.23 ;
      RECT 2.215 0.35 2.315 1.23 ;
      RECT 0.785 1.05 1.505 1.14 ;
      RECT 1.415 0.25 1.505 1.14 ;
      RECT 2.2 0.89 2.315 1.23 ;
      RECT 1.775 0.89 1.865 1.23 ;
      RECT 1.415 0.89 1.865 0.98 ;
      RECT 2.175 0.35 2.315 0.44 ;
      RECT 0.865 0.25 1.505 0.34 ;
      RECT 0.045 1.05 0.185 1.14 ;
      RECT 0.045 0.25 0.135 1.14 ;
      RECT 0.945 0.795 1.325 0.885 ;
      RECT 0.945 0.495 1.035 0.885 ;
      RECT 0.685 0.495 1.035 0.585 ;
      RECT 0.685 0.265 0.775 0.585 ;
      RECT 0.045 0.265 0.775 0.355 ;
      RECT 0.045 0.25 0.185 0.355 ;
  END
END SDFFSX2H7R

MACRO SDFFTRQX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFTRQX0P5H7R 0 0 ;
  SIZE 6.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.8 1.48 ;
        RECT 6.38 1.005 6.47 1.48 ;
        RECT 5.87 1.05 5.96 1.48 ;
        RECT 4.74 1.125 4.91 1.48 ;
        RECT 3.35 1.005 3.44 1.48 ;
        RECT 2.23 1.185 2.32 1.48 ;
        RECT 1.78 1.07 1.87 1.48 ;
        RECT 0.34 1.07 0.43 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.8 0.08 ;
        RECT 6.38 -0.08 6.47 0.375 ;
        RECT 5.805 -0.08 5.955 0.175 ;
        RECT 4.585 -0.08 4.735 0.175 ;
        RECT 3.025 -0.08 3.175 0.175 ;
        RECT 1.945 -0.08 2.035 0.33 ;
        RECT 0.34 -0.08 0.43 0.33 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 5.645 0.54 5.76 0.775 ;
      LAYER MET2 ;
        RECT 5.65 0.425 5.75 0.96 ;
      LAYER VIA1 ;
        RECT 5.655 0.655 5.745 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.855 0.6 1.995 0.795 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.63 0.225 6.745 1.045 ;
      LAYER MET2 ;
        RECT 6.65 0.18 6.75 0.56 ;
      LAYER VIA1 ;
        RECT 6.655 0.255 6.745 0.345 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.4 0.6 1.545 0.79 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.86 1.14 1.045 1.23 ;
        RECT 0.86 0.465 0.95 1.23 ;
        RECT 0.225 0.465 0.95 0.555 ;
        RECT 0.225 0.44 0.375 0.555 ;
        RECT 0.225 0.44 0.34 0.58 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 0.655 0.59 0.8 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 6.15 0.27 6.24 1.05 ;
      RECT 4.43 0.485 4.75 0.575 ;
      RECT 4.66 0.363 4.75 0.575 ;
      RECT 5.841 0.385 6.24 0.475 ;
      RECT 5.802 0.327 5.841 0.456 ;
      RECT 5.756 0.285 5.802 0.413 ;
      RECT 5.756 0.366 5.879 0.413 ;
      RECT 5.71 0.239 5.756 0.367 ;
      RECT 4.706 0.318 4.796 0.401 ;
      RECT 5.664 0.193 5.71 0.321 ;
      RECT 4.75 0.273 4.842 0.355 ;
      RECT 5.626 0.239 5.756 0.279 ;
      RECT 4.796 0.227 4.914 0.279 ;
      RECT 4.842 0.187 4.876 0.315 ;
      RECT 4.876 0.17 5.664 0.26 ;
      RECT 5 1.14 5.72 1.23 ;
      RECT 5.63 0.87 5.72 1.23 ;
      RECT 5 0.945 5.09 1.23 ;
      RECT 4.07 0.96 4.6 1.05 ;
      RECT 4.51 0.945 5.09 1.035 ;
      RECT 5.63 0.87 6.06 0.96 ;
      RECT 5.97 0.615 6.06 0.96 ;
      RECT 4.07 0.35 4.16 1.05 ;
      RECT 3.99 0.35 4.16 0.465 ;
      RECT 5.445 0.36 5.535 1.05 ;
      RECT 5.08 0.585 5.535 0.675 ;
      RECT 5.445 0.36 5.595 0.45 ;
      RECT 5.18 0.765 5.27 1.05 ;
      RECT 4.9 0.765 5.27 0.855 ;
      RECT 4.25 0.665 4.38 0.83 ;
      RECT 4.9 0.405 4.99 0.855 ;
      RECT 4.25 0.665 4.99 0.755 ;
      RECT 4.25 0.17 4.34 0.83 ;
      RECT 2.7 0.285 2.79 0.605 ;
      RECT 3.805 0.17 3.895 0.58 ;
      RECT 4.9 0.405 5.245 0.495 ;
      RECT 5.155 0.35 5.295 0.44 ;
      RECT 2.7 0.285 3.355 0.375 ;
      RECT 3.265 0.17 3.355 0.375 ;
      RECT 3.265 0.17 4.34 0.26 ;
      RECT 3.53 1.14 3.98 1.23 ;
      RECT 3.89 0.715 3.98 1.23 ;
      RECT 2.49 1.14 3.195 1.23 ;
      RECT 3.105 0.825 3.195 1.23 ;
      RECT 3.53 0.825 3.62 1.23 ;
      RECT 2.49 0.915 2.58 1.23 ;
      RECT 2.34 0.915 2.58 1.005 ;
      RECT 3.105 0.825 3.62 0.915 ;
      RECT 2.34 0.465 2.43 1.005 ;
      RECT 3.71 0.721 3.8 1.05 ;
      RECT 3.686 0.721 3.8 0.767 ;
      RECT 3.64 0.465 3.715 0.732 ;
      RECT 3.64 0.679 3.761 0.732 ;
      RECT 3.625 0.35 3.64 0.702 ;
      RECT 2.945 0.465 3.715 0.555 ;
      RECT 3.5 0.35 3.64 0.555 ;
      RECT 2.8 0.695 2.89 1.025 ;
      RECT 2.52 0.695 2.97 0.785 ;
      RECT 2.88 0.645 3.535 0.735 ;
      RECT 2.52 0.225 2.61 0.785 ;
      RECT 2.425 0.225 2.61 0.315 ;
      RECT 1.04 0.17 1.13 1.05 ;
      RECT 2.11 0.42 2.2 0.615 ;
      RECT 1.495 0.42 2.2 0.51 ;
      RECT 1.495 0.17 1.585 0.51 ;
      RECT 0.785 0.25 1.13 0.34 ;
      RECT 1.04 0.17 1.585 0.26 ;
      RECT 2.05 0.89 2.14 1.065 ;
      RECT 1.31 0.89 1.4 1.06 ;
      RECT 1.22 0.89 2.14 0.98 ;
      RECT 1.22 0.35 1.31 0.98 ;
      RECT 1.22 0.35 1.36 0.455 ;
      RECT 0.045 0.89 0.16 1.065 ;
      RECT 0.045 0.89 0.77 0.98 ;
      RECT 0.68 0.7 0.77 0.98 ;
      RECT 0.045 0.26 0.135 1.065 ;
      RECT 0.045 0.26 0.185 0.35 ;
  END
END SDFFTRQX0P5H7R

MACRO SDFFTRQX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFTRQX1H7R 0 0 ;
  SIZE 6.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 6.8 1.48 ;
        RECT 6.255 1.05 6.345 1.48 ;
        RECT 5.245 1.095 5.385 1.48 ;
        RECT 3.915 1.225 4.055 1.48 ;
        RECT 2.65 1.12 2.79 1.48 ;
        RECT 1.48 1.225 1.62 1.48 ;
        RECT 0.315 1.075 0.455 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 6.8 0.08 ;
        RECT 6.04 -0.08 6.13 0.33 ;
        RECT 5.19 -0.08 5.33 0.285 ;
        RECT 3.805 -0.08 3.945 0.16 ;
        RECT 2.74 -0.08 2.88 0.175 ;
        RECT 2.22 -0.08 2.36 0.16 ;
        RECT 0.34 -0.08 0.43 0.33 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 2.425 0.455 2.685 0.615 ;
      LAYER MET2 ;
        RECT 2.45 0.225 2.55 0.76 ;
      LAYER VIA1 ;
        RECT 2.455 0.455 2.545 0.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.835 0.54 1.95 0.775 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.525 0.655 6.615 0.985 ;
        RECT 6.425 0.655 6.615 0.745 ;
        RECT 6.425 0.24 6.515 0.745 ;
      LAYER MET2 ;
        RECT 6.45 0.425 6.55 0.96 ;
      LAYER VIA1 ;
        RECT 6.455 0.655 6.545 0.745 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.365 0.625 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.755 0.455 0.895 0.565 ;
        RECT 0.225 0.455 0.895 0.545 ;
        RECT 0.225 0.455 0.315 0.605 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.415 0.635 0.595 0.785 ;
      LAYER MET2 ;
        RECT 0.45 0.415 0.55 0.945 ;
      LAYER VIA1 ;
        RECT 0.455 0.64 0.545 0.73 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.586 1.075 6.165 1.165 ;
      RECT 6.075 0.555 6.165 1.165 ;
      RECT 5.556 1.022 5.586 1.15 ;
      RECT 5.51 0.984 5.556 1.112 ;
      RECT 5.51 1.056 5.624 1.112 ;
      RECT 5.464 0.938 5.51 1.066 ;
      RECT 5.426 0.915 5.464 1.024 ;
      RECT 4.555 0.915 5.464 1.005 ;
      RECT 4.555 0.35 4.645 1.005 ;
      RECT 4.44 0.35 4.645 0.44 ;
      RECT 5.895 0.555 5.985 0.985 ;
      RECT 5.075 0.555 5.985 0.645 ;
      RECT 5.77 0.275 5.86 0.645 ;
      RECT 5.65 0.735 5.74 0.97 ;
      RECT 4.78 0.735 5.74 0.825 ;
      RECT 4.78 0.715 4.93 0.825 ;
      RECT 4.78 0.17 4.87 0.825 ;
      RECT 4.78 0.375 5.63 0.465 ;
      RECT 5.54 0.24 5.63 0.465 ;
      RECT 3.55 0.28 4.004 0.37 ;
      RECT 3.55 0.28 4.05 0.347 ;
      RECT 3.966 0.261 4.076 0.311 ;
      RECT 3.55 0.17 3.64 0.37 ;
      RECT 4.004 0.219 4.114 0.279 ;
      RECT 4.05 0.183 4.076 0.311 ;
      RECT 4.076 0.17 4.87 0.26 ;
      RECT 3.415 0.17 3.64 0.26 ;
      RECT 4.24 1.14 4.785 1.23 ;
      RECT 3.11 1.14 3.78 1.23 ;
      RECT 3.69 1.045 3.78 1.23 ;
      RECT 4.24 1.045 4.33 1.23 ;
      RECT 3.11 0.524 3.2 1.23 ;
      RECT 3.69 1.045 4.33 1.135 ;
      RECT 2.4 0.94 2.49 1.08 ;
      RECT 2.4 0.94 3.2 1.03 ;
      RECT 3.085 0.443 3.11 0.572 ;
      RECT 3.041 0.479 3.156 0.537 ;
      RECT 2.995 0.275 3.085 0.492 ;
      RECT 2.465 0.275 3.085 0.365 ;
      RECT 3.84 0.865 4.335 0.955 ;
      RECT 4.245 0.35 4.335 0.955 ;
      RECT 3.84 0.72 3.93 0.955 ;
      RECT 3.77 0.72 3.93 0.81 ;
      RECT 4.155 0.35 4.335 0.44 ;
      RECT 3.455 0.54 3.545 1.045 ;
      RECT 4.055 0.54 4.145 0.69 ;
      RECT 3.29 0.54 4.145 0.63 ;
      RECT 3.29 0.35 3.38 0.63 ;
      RECT 3.225 0.35 3.38 0.44 ;
      RECT 0.795 1.055 1.125 1.145 ;
      RECT 2.22 0.358 2.31 1.135 ;
      RECT 1.035 1.045 2.31 1.135 ;
      RECT 2.22 0.76 2.94 0.85 ;
      RECT 2.85 0.675 2.94 0.85 ;
      RECT 2.192 0.276 2.22 0.404 ;
      RECT 2.146 0.239 2.192 0.367 ;
      RECT 2.146 0.313 2.266 0.367 ;
      RECT 0.92 0.17 1.01 0.33 ;
      RECT 2.1 0.193 2.146 0.321 ;
      RECT 2.062 0.17 2.1 0.279 ;
      RECT 0.92 0.17 2.1 0.26 ;
      RECT 1.135 0.865 2.13 0.955 ;
      RECT 2.04 0.434 2.13 0.955 ;
      RECT 2.024 0.358 2.04 0.486 ;
      RECT 1.986 0.434 2.13 0.459 ;
      RECT 1.245 0.35 2.024 0.44 ;
      RECT 1.245 0.389 2.086 0.44 ;
      RECT 0.045 0.875 0.8 0.965 ;
      RECT 0.71 0.655 0.8 0.965 ;
      RECT 0.045 0.28 0.135 0.965 ;
      RECT 0.71 0.655 1.25 0.745 ;
      RECT 1.16 0.53 1.25 0.745 ;
      RECT 0.045 0.28 0.185 0.37 ;
  END
END SDFFTRQX1H7R

MACRO SDFFTRQX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFTRQX2H7R 0 0 ;
  SIZE 7 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7 1.48 ;
        RECT 6.795 0.995 6.885 1.48 ;
        RECT 6.255 0.995 6.345 1.48 ;
        RECT 5.245 1.095 5.385 1.48 ;
        RECT 3.915 1.225 4.055 1.48 ;
        RECT 2.65 1.075 2.79 1.48 ;
        RECT 1.48 1.225 1.62 1.48 ;
        RECT 0.315 1.075 0.455 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7 0.08 ;
        RECT 6.715 -0.08 6.805 0.385 ;
        RECT 6.04 -0.08 6.13 0.33 ;
        RECT 5.19 -0.08 5.33 0.285 ;
        RECT 3.805 -0.08 3.945 0.16 ;
        RECT 2.74 -0.08 2.88 0.175 ;
        RECT 2.22 -0.08 2.36 0.16 ;
        RECT 0.34 -0.08 0.43 0.33 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 2.545 0.455 2.775 0.545 ;
        RECT 2.545 0.455 2.685 0.615 ;
      LAYER MET2 ;
        RECT 2.65 0.23 2.75 0.76 ;
      LAYER VIA1 ;
        RECT 2.655 0.455 2.745 0.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.835 0.54 1.95 0.775 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.525 0.655 6.615 1.105 ;
        RECT 6.425 0.655 6.615 0.745 ;
        RECT 6.425 0.24 6.515 0.745 ;
      LAYER MET2 ;
        RECT 6.45 0.425 6.55 0.96 ;
      LAYER VIA1 ;
        RECT 6.455 0.655 6.545 0.745 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.365 0.625 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.755 0.455 0.895 0.565 ;
        RECT 0.225 0.455 0.895 0.545 ;
        RECT 0.225 0.455 0.315 0.645 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.415 0.65 0.595 0.8 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.586 1.075 6.165 1.165 ;
      RECT 6.075 0.555 6.165 1.165 ;
      RECT 5.556 1.022 5.586 1.15 ;
      RECT 5.51 0.984 5.556 1.112 ;
      RECT 5.51 1.056 5.624 1.112 ;
      RECT 5.464 0.938 5.51 1.066 ;
      RECT 5.426 0.915 5.464 1.024 ;
      RECT 4.52 0.915 5.464 1.005 ;
      RECT 4.52 0.35 4.61 1.005 ;
      RECT 4.435 0.35 4.61 0.44 ;
      RECT 5.895 0.555 5.985 0.985 ;
      RECT 5.075 0.555 5.985 0.645 ;
      RECT 5.77 0.295 5.86 0.645 ;
      RECT 5.65 0.735 5.74 0.97 ;
      RECT 4.78 0.735 5.74 0.825 ;
      RECT 4.78 0.715 4.93 0.825 ;
      RECT 4.78 0.17 4.87 0.825 ;
      RECT 4.78 0.375 5.63 0.465 ;
      RECT 5.54 0.295 5.63 0.465 ;
      RECT 3.55 0.28 4.004 0.37 ;
      RECT 3.55 0.28 4.05 0.347 ;
      RECT 3.966 0.261 4.076 0.311 ;
      RECT 3.55 0.17 3.64 0.37 ;
      RECT 4.004 0.219 4.114 0.279 ;
      RECT 4.05 0.183 4.076 0.311 ;
      RECT 4.076 0.17 4.87 0.26 ;
      RECT 3.415 0.17 3.64 0.26 ;
      RECT 4.24 1.14 4.785 1.23 ;
      RECT 3.11 1.14 3.78 1.23 ;
      RECT 3.69 1.045 3.78 1.23 ;
      RECT 4.24 1.045 4.33 1.23 ;
      RECT 3.11 0.524 3.2 1.23 ;
      RECT 3.69 1.045 4.33 1.135 ;
      RECT 2.4 0.885 2.49 1.025 ;
      RECT 2.4 0.885 3.2 0.975 ;
      RECT 3.085 0.443 3.11 0.572 ;
      RECT 3.041 0.479 3.156 0.537 ;
      RECT 2.995 0.275 3.085 0.492 ;
      RECT 2.465 0.275 3.085 0.365 ;
      RECT 3.84 0.865 4.33 0.955 ;
      RECT 4.24 0.35 4.33 0.955 ;
      RECT 3.84 0.72 3.93 0.955 ;
      RECT 3.77 0.72 3.93 0.81 ;
      RECT 4.155 0.35 4.33 0.44 ;
      RECT 3.455 0.54 3.545 1.045 ;
      RECT 4.055 0.54 4.145 0.69 ;
      RECT 3.29 0.54 4.145 0.63 ;
      RECT 3.29 0.35 3.38 0.63 ;
      RECT 3.225 0.35 3.38 0.44 ;
      RECT 0.795 1.07 1.125 1.16 ;
      RECT 2.22 0.358 2.31 1.135 ;
      RECT 1.035 1.045 2.31 1.135 ;
      RECT 2.22 0.705 2.965 0.795 ;
      RECT 2.825 0.685 2.965 0.795 ;
      RECT 2.192 0.276 2.22 0.404 ;
      RECT 2.146 0.239 2.192 0.367 ;
      RECT 2.146 0.313 2.266 0.367 ;
      RECT 0.92 0.17 1.01 0.33 ;
      RECT 2.1 0.193 2.146 0.321 ;
      RECT 2.062 0.17 2.1 0.279 ;
      RECT 0.92 0.17 2.1 0.26 ;
      RECT 1.135 0.865 2.13 0.955 ;
      RECT 2.04 0.434 2.13 0.955 ;
      RECT 2.024 0.358 2.04 0.486 ;
      RECT 1.986 0.434 2.13 0.459 ;
      RECT 1.245 0.35 2.024 0.44 ;
      RECT 1.245 0.389 2.086 0.44 ;
      RECT 0.045 0.89 0.8 0.98 ;
      RECT 0.71 0.655 0.8 0.98 ;
      RECT 0.045 0.28 0.135 0.98 ;
      RECT 0.71 0.655 1.25 0.745 ;
      RECT 1.16 0.53 1.25 0.745 ;
      RECT 0.045 0.28 0.185 0.37 ;
  END
END SDFFTRQX2H7R

MACRO SDFFTRQX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFTRQX3H7R 0 0 ;
  SIZE 7 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7 1.48 ;
        RECT 6.795 0.995 6.885 1.48 ;
        RECT 6.255 0.995 6.345 1.48 ;
        RECT 5.245 1.095 5.385 1.48 ;
        RECT 3.915 1.225 4.055 1.48 ;
        RECT 2.65 1.225 2.79 1.48 ;
        RECT 1.48 1.225 1.62 1.48 ;
        RECT 0.34 1.07 0.43 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7 0.08 ;
        RECT 6.715 -0.08 6.805 0.385 ;
        RECT 6.04 -0.08 6.13 0.38 ;
        RECT 5.19 -0.08 5.33 0.285 ;
        RECT 3.805 -0.08 3.945 0.16 ;
        RECT 2.74 -0.08 2.88 0.175 ;
        RECT 2.22 -0.08 2.36 0.16 ;
        RECT 0.34 -0.08 0.43 0.335 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 2.42 0.455 2.685 0.615 ;
      LAYER MET2 ;
        RECT 2.45 0.225 2.55 0.76 ;
      LAYER VIA1 ;
        RECT 2.455 0.455 2.545 0.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.835 0.54 1.95 0.775 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.525 0.655 6.615 0.97 ;
        RECT 6.425 0.655 6.615 0.745 ;
        RECT 6.425 0.24 6.515 0.745 ;
      LAYER MET2 ;
        RECT 6.45 0.425 6.55 0.96 ;
      LAYER VIA1 ;
        RECT 6.455 0.655 6.545 0.745 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.365 0.625 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END RN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.755 0.455 0.895 0.565 ;
        RECT 0.225 0.455 0.895 0.545 ;
        RECT 0.225 0.455 0.315 0.645 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.415 0.65 0.595 0.8 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.586 1.075 6.165 1.165 ;
      RECT 6.075 0.555 6.165 1.165 ;
      RECT 5.556 1.022 5.586 1.15 ;
      RECT 5.51 0.984 5.556 1.112 ;
      RECT 5.51 1.056 5.624 1.112 ;
      RECT 5.464 0.938 5.51 1.066 ;
      RECT 5.426 0.915 5.464 1.024 ;
      RECT 4.52 0.915 5.464 1.005 ;
      RECT 4.52 0.35 4.61 1.005 ;
      RECT 4.435 0.35 4.61 0.465 ;
      RECT 5.895 0.555 5.985 0.985 ;
      RECT 5.075 0.555 5.985 0.645 ;
      RECT 5.77 0.24 5.86 0.645 ;
      RECT 5.65 0.735 5.74 0.97 ;
      RECT 4.78 0.735 5.74 0.825 ;
      RECT 4.78 0.715 4.93 0.825 ;
      RECT 4.78 0.17 4.87 0.825 ;
      RECT 4.78 0.375 5.63 0.465 ;
      RECT 5.54 0.24 5.63 0.465 ;
      RECT 3.55 0.28 4.004 0.37 ;
      RECT 3.55 0.28 4.05 0.347 ;
      RECT 3.966 0.261 4.076 0.311 ;
      RECT 3.55 0.17 3.64 0.37 ;
      RECT 4.004 0.219 4.114 0.279 ;
      RECT 4.05 0.183 4.076 0.311 ;
      RECT 4.076 0.17 4.87 0.26 ;
      RECT 3.415 0.17 3.64 0.26 ;
      RECT 4.24 1.14 4.785 1.23 ;
      RECT 3.11 1.14 3.78 1.23 ;
      RECT 3.69 1.045 3.78 1.23 ;
      RECT 2.4 1.02 2.49 1.16 ;
      RECT 4.24 1.045 4.33 1.23 ;
      RECT 3.11 0.524 3.2 1.23 ;
      RECT 3.69 1.045 4.33 1.135 ;
      RECT 2.4 1.045 3.2 1.135 ;
      RECT 3.085 0.443 3.11 0.572 ;
      RECT 3.041 0.479 3.156 0.537 ;
      RECT 2.995 0.275 3.085 0.492 ;
      RECT 2.465 0.275 3.085 0.365 ;
      RECT 3.84 0.865 4.33 0.955 ;
      RECT 4.24 0.35 4.33 0.955 ;
      RECT 3.84 0.72 3.93 0.955 ;
      RECT 3.77 0.72 3.93 0.81 ;
      RECT 4.155 0.35 4.33 0.44 ;
      RECT 3.455 0.54 3.545 1.045 ;
      RECT 4.055 0.54 4.145 0.69 ;
      RECT 3.29 0.54 4.145 0.63 ;
      RECT 3.29 0.35 3.38 0.63 ;
      RECT 3.225 0.35 3.38 0.44 ;
      RECT 0.795 1.07 1.125 1.16 ;
      RECT 2.22 0.358 2.31 1.135 ;
      RECT 1.035 1.045 2.31 1.135 ;
      RECT 2.22 0.76 2.94 0.85 ;
      RECT 2.85 0.615 2.94 0.85 ;
      RECT 2.192 0.276 2.22 0.404 ;
      RECT 2.146 0.239 2.192 0.367 ;
      RECT 0.92 0.17 1.01 0.36 ;
      RECT 2.146 0.313 2.266 0.367 ;
      RECT 2.1 0.193 2.146 0.321 ;
      RECT 2.062 0.17 2.1 0.279 ;
      RECT 0.92 0.17 2.1 0.26 ;
      RECT 1.135 0.865 2.13 0.955 ;
      RECT 2.04 0.434 2.13 0.955 ;
      RECT 2.024 0.358 2.04 0.486 ;
      RECT 1.986 0.434 2.13 0.459 ;
      RECT 1.245 0.35 2.024 0.44 ;
      RECT 1.245 0.389 2.086 0.44 ;
      RECT 0.045 0.89 0.8 0.98 ;
      RECT 0.71 0.655 0.8 0.98 ;
      RECT 0.045 0.28 0.135 0.98 ;
      RECT 0.71 0.655 1.25 0.745 ;
      RECT 1.16 0.53 1.25 0.745 ;
      RECT 0.045 0.28 0.185 0.37 ;
  END
END SDFFTRQX3H7R

MACRO SDFFX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFX0P5H7R 0 0 ;
  SIZE 7 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7 1.48 ;
        RECT 6.32 0.995 6.41 1.48 ;
        RECT 5.76 1.01 5.85 1.48 ;
        RECT 4.75 1.105 4.89 1.48 ;
        RECT 3.54 1.24 3.68 1.48 ;
        RECT 2.67 1.24 2.81 1.48 ;
        RECT 1.215 1.24 1.355 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7 0.08 ;
        RECT 6.435 -0.08 6.525 0.345 ;
        RECT 5.715 -0.08 5.805 0.33 ;
        RECT 4.76 -0.08 4.9 0.275 ;
        RECT 3.54 -0.08 3.68 0.16 ;
        RECT 2.64 -0.08 2.73 0.235 ;
        RECT 1.025 -0.08 1.165 0.16 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.21 0.65 3.48 0.75 ;
      LAYER MET2 ;
        RECT 3.25 0.43 3.35 0.96 ;
      LAYER VIA1 ;
        RECT 3.255 0.655 3.345 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.27 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.005 0.825 6.165 0.98 ;
        RECT 6.075 0.35 6.165 0.98 ;
      LAYER MET2 ;
        RECT 6.05 0.63 6.15 1.16 ;
      LAYER VIA1 ;
        RECT 6.055 0.855 6.145 0.945 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.545 0.825 6.775 0.975 ;
        RECT 6.685 0.255 6.775 0.975 ;
      LAYER MET2 ;
        RECT 6.65 0.625 6.75 1.16 ;
      LAYER VIA1 ;
        RECT 6.655 0.855 6.745 0.945 ;
    END
  END QN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.34 0.508 1.43 0.67 ;
        RECT 0.655 0.468 1.395 0.535 ;
        RECT 0.655 0.445 1.349 0.535 ;
        RECT 1.311 0.508 1.43 0.55 ;
        RECT 0.655 0.445 0.775 0.6 ;
        RECT 0.655 0.445 0.745 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.015 0.625 1.19 0.79 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.4 0.255 5.49 1.005 ;
      RECT 4.81 0.56 5.49 0.65 ;
      RECT 6.255 0.49 6.595 0.58 ;
      RECT 5.4 0.455 5.985 0.545 ;
      RECT 5.895 0.17 5.985 0.545 ;
      RECT 6.255 0.17 6.345 0.58 ;
      RECT 5.895 0.17 6.345 0.26 ;
      RECT 4.99 1.135 5.67 1.225 ;
      RECT 5.58 0.645 5.67 1.225 ;
      RECT 4.99 0.925 5.08 1.225 ;
      RECT 4.04 0.925 5.08 1.015 ;
      RECT 4.04 0.35 4.185 1.015 ;
      RECT 5.58 0.645 5.955 0.735 ;
      RECT 5.17 0.74 5.26 1.045 ;
      RECT 4.275 0.74 5.26 0.83 ;
      RECT 4.275 0.17 4.365 0.83 ;
      RECT 2.275 0.325 2.365 0.575 ;
      RECT 4.275 0.365 5.26 0.455 ;
      RECT 5.17 0.305 5.26 0.455 ;
      RECT 2.275 0.325 2.94 0.415 ;
      RECT 2.85 0.17 2.94 0.415 ;
      RECT 3.275 0.25 3.885 0.34 ;
      RECT 3.795 0.17 4.365 0.26 ;
      RECT 2.85 0.17 3.365 0.26 ;
      RECT 3.825 1.14 4.265 1.23 ;
      RECT 1.915 1.125 2.48 1.215 ;
      RECT 3.825 0.43 3.915 1.23 ;
      RECT 2.39 1.045 3.915 1.135 ;
      RECT 1.915 0.48 2.005 1.215 ;
      RECT 3.26 0.43 3.915 0.52 ;
      RECT 3 0.865 3.735 0.955 ;
      RECT 3.645 0.635 3.735 0.955 ;
      RECT 3.03 0.35 3.12 0.955 ;
      RECT 2.515 0.505 3.12 0.595 ;
      RECT 2.095 0.24 2.185 1.01 ;
      RECT 2.095 0.725 2.89 0.815 ;
      RECT 1.685 1.06 1.825 1.23 ;
      RECT 1.735 0.17 1.825 1.23 ;
      RECT 0.705 1.06 1.825 1.15 ;
      RECT 1.735 0.17 1.88 0.375 ;
      RECT 0.505 0.25 1.35 0.34 ;
      RECT 1.26 0.17 1.88 0.26 ;
      RECT 0.4 0.88 1.645 0.97 ;
      RECT 1.555 0.35 1.645 0.97 ;
      RECT 0.835 0.725 0.925 0.97 ;
      RECT 0.4 0.505 0.49 0.97 ;
      RECT 1.505 0.35 1.645 0.44 ;
  END
END SDFFX0P5H7R

MACRO SDFFX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFX1H7R 0 0 ;
  SIZE 7 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7 1.48 ;
        RECT 6.315 0.87 6.405 1.48 ;
        RECT 5.76 1.07 5.85 1.48 ;
        RECT 4.73 1.09 4.87 1.48 ;
        RECT 3.54 1.24 3.68 1.48 ;
        RECT 2.67 1.24 2.81 1.48 ;
        RECT 1.2 1.24 1.34 1.48 ;
        RECT 0.07 1.015 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7 0.08 ;
        RECT 6.465 -0.08 6.555 0.345 ;
        RECT 5.695 -0.08 5.785 0.365 ;
        RECT 4.82 -0.08 4.96 0.275 ;
        RECT 3.54 -0.08 3.68 0.16 ;
        RECT 2.64 -0.08 2.73 0.185 ;
        RECT 1.025 -0.08 1.165 0.16 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.335 0.61 3.575 0.75 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.055 0.35 6.195 1.19 ;
      LAYER MET2 ;
        RECT 6.05 0.84 6.15 1.22 ;
      LAYER VIA1 ;
        RECT 6.055 1.055 6.145 1.145 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.585 0.855 6.815 0.945 ;
        RECT 6.725 0.245 6.815 0.945 ;
        RECT 6.585 0.855 6.675 1.195 ;
      LAYER MET2 ;
        RECT 6.65 0.625 6.75 1.16 ;
      LAYER VIA1 ;
        RECT 6.655 0.855 6.745 0.945 ;
    END
  END QN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.325 0.43 1.415 0.625 ;
        RECT 0.655 0.43 1.415 0.52 ;
        RECT 0.655 0.43 0.745 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.045 0.61 1.195 0.79 ;
      LAYER MET2 ;
        RECT 1.04 0.425 1.14 0.96 ;
      LAYER VIA1 ;
        RECT 1.045 0.655 1.135 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.4 0.545 5.49 1.005 ;
      RECT 6.285 0.56 6.62 0.65 ;
      RECT 4.81 0.545 5.49 0.635 ;
      RECT 5.875 0.17 5.965 0.615 ;
      RECT 6.285 0.17 6.375 0.65 ;
      RECT 5.425 0.525 5.965 0.615 ;
      RECT 5.425 0.31 5.515 0.615 ;
      RECT 5.875 0.17 6.375 0.26 ;
      RECT 4.97 1.14 5.67 1.23 ;
      RECT 5.58 0.705 5.67 1.23 ;
      RECT 4.97 0.91 5.06 1.23 ;
      RECT 4.04 0.91 5.06 1 ;
      RECT 4.04 0.35 4.13 1 ;
      RECT 5.58 0.705 5.74 0.795 ;
      RECT 4.04 0.35 4.185 0.44 ;
      RECT 5.155 0.73 5.245 1.045 ;
      RECT 4.275 0.73 5.245 0.82 ;
      RECT 4.275 0.17 4.365 0.82 ;
      RECT 2.275 0.275 2.365 0.575 ;
      RECT 4.275 0.365 5.285 0.455 ;
      RECT 5.195 0.275 5.285 0.455 ;
      RECT 2.275 0.275 2.91 0.365 ;
      RECT 2.82 0.17 2.91 0.365 ;
      RECT 3.36 0.25 3.86 0.34 ;
      RECT 3.77 0.17 4.365 0.26 ;
      RECT 2.82 0.17 3.45 0.26 ;
      RECT 3.825 1.14 4.265 1.23 ;
      RECT 1.915 1.125 2.48 1.215 ;
      RECT 3.825 1.045 3.95 1.23 ;
      RECT 3.86 0.43 3.95 1.23 ;
      RECT 2.39 1.045 3.95 1.135 ;
      RECT 1.915 0.48 2.005 1.215 ;
      RECT 3.25 1.02 3.39 1.135 ;
      RECT 3.26 0.43 3.95 0.52 ;
      RECT 3.005 0.35 3.145 0.955 ;
      RECT 3.005 0.84 3.77 0.93 ;
      RECT 3.68 0.665 3.77 0.93 ;
      RECT 2.515 0.475 3.145 0.565 ;
      RECT 3 0.35 3.145 0.565 ;
      RECT 2.095 0.24 2.185 1.035 ;
      RECT 2.095 0.8 2.915 0.89 ;
      RECT 2.825 0.675 2.915 0.89 ;
      RECT 0.705 1.06 1.825 1.15 ;
      RECT 1.735 0.17 1.825 1.15 ;
      RECT 1.735 0.17 1.88 0.365 ;
      RECT 0.505 0.25 1.35 0.34 ;
      RECT 1.26 0.17 1.88 0.26 ;
      RECT 0.4 0.88 1.645 0.97 ;
      RECT 1.505 0.35 1.645 0.97 ;
      RECT 0.865 0.725 0.955 0.97 ;
      RECT 0.4 0.505 0.49 0.97 ;
  END
END SDFFX1H7R

MACRO SDFFX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFX2H7R 0 0 ;
  SIZE 7.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7.2 1.48 ;
        RECT 6.925 1.055 7.015 1.48 ;
        RECT 6.395 1.07 6.485 1.48 ;
        RECT 5.855 1.07 5.945 1.48 ;
        RECT 4.84 1.09 4.98 1.48 ;
        RECT 3.57 1.24 3.71 1.48 ;
        RECT 2.7 1.24 2.84 1.48 ;
        RECT 1.215 1.24 1.355 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7.2 0.08 ;
        RECT 6.935 -0.08 7.025 0.33 ;
        RECT 6.395 -0.08 6.485 0.33 ;
        RECT 5.855 -0.08 5.945 0.33 ;
        RECT 4.85 -0.08 4.99 0.275 ;
        RECT 3.57 -0.08 3.71 0.16 ;
        RECT 2.67 -0.08 2.76 0.185 ;
        RECT 1.025 -0.08 1.165 0.16 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.35 0.655 3.575 0.775 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.125 0.805 6.545 0.895 ;
        RECT 6.455 0.435 6.545 0.895 ;
        RECT 6.215 0.435 6.545 0.525 ;
        RECT 6.215 0.235 6.305 0.525 ;
        RECT 6.125 0.805 6.215 1.17 ;
        RECT 6.1 0.235 6.305 0.325 ;
      LAYER MET2 ;
        RECT 6.45 0.425 6.55 0.96 ;
      LAYER VIA1 ;
        RECT 6.455 0.655 6.545 0.745 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.655 0.21 6.745 1.13 ;
      LAYER MET2 ;
        RECT 6.65 0.625 6.75 1.16 ;
      LAYER VIA1 ;
        RECT 6.655 0.855 6.745 0.945 ;
    END
  END QN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.34 0.445 1.43 0.72 ;
        RECT 0.655 0.445 1.43 0.535 ;
        RECT 0.655 0.445 0.745 0.775 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.055 0.625 1.235 0.775 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.495 0.545 5.585 1.005 ;
      RECT 6.025 0.625 6.34 0.715 ;
      RECT 4.85 0.545 5.585 0.635 ;
      RECT 6.025 0.525 6.115 0.715 ;
      RECT 5.525 0.525 6.115 0.615 ;
      RECT 5.525 0.32 5.615 0.615 ;
      RECT 5.525 0.32 5.7 0.41 ;
      RECT 5.07 1.095 5.765 1.185 ;
      RECT 5.675 0.705 5.765 1.185 ;
      RECT 5.07 0.91 5.16 1.185 ;
      RECT 4.07 0.91 5.16 1 ;
      RECT 4.07 0.885 4.21 1 ;
      RECT 4.07 0.35 4.16 1 ;
      RECT 5.675 0.705 5.89 0.795 ;
      RECT 4.07 0.35 4.215 0.44 ;
      RECT 5.25 0.73 5.34 1.005 ;
      RECT 4.305 0.73 5.34 0.82 ;
      RECT 4.305 0.17 4.395 0.82 ;
      RECT 2.305 0.275 2.395 0.575 ;
      RECT 4.305 0.365 5.335 0.455 ;
      RECT 5.245 0.295 5.335 0.455 ;
      RECT 2.305 0.275 2.94 0.365 ;
      RECT 2.85 0.17 2.94 0.365 ;
      RECT 3.491 0.25 3.915 0.34 ;
      RECT 3.449 0.191 3.491 0.319 ;
      RECT 3.411 0.25 3.915 0.279 ;
      RECT 3.825 0.17 4.395 0.26 ;
      RECT 2.85 0.231 3.529 0.26 ;
      RECT 2.85 0.17 3.449 0.26 ;
      RECT 3.89 1.14 4.295 1.23 ;
      RECT 1.945 1.125 2.51 1.215 ;
      RECT 2.42 1.06 3.98 1.15 ;
      RECT 1.945 0.48 2.035 1.215 ;
      RECT 3.89 0.43 3.98 1.23 ;
      RECT 3.29 0.43 3.98 0.52 ;
      RECT 3.29 0.415 3.43 0.52 ;
      RECT 3.035 0.88 3.765 0.97 ;
      RECT 3.675 0.66 3.765 0.97 ;
      RECT 3.035 0.35 3.175 0.97 ;
      RECT 2.545 0.475 3.175 0.565 ;
      RECT 2.125 0.225 2.215 1.03 ;
      RECT 2.125 0.8 2.945 0.89 ;
      RECT 2.855 0.66 2.945 0.89 ;
      RECT 0.715 1.06 1.855 1.15 ;
      RECT 1.765 0.17 1.855 1.15 ;
      RECT 1.765 0.17 1.91 0.365 ;
      RECT 0.525 0.25 1.35 0.34 ;
      RECT 1.26 0.17 1.91 0.26 ;
      RECT 0.4 0.88 1.675 0.97 ;
      RECT 1.535 0.35 1.675 0.97 ;
      RECT 0.87 0.725 0.96 0.97 ;
      RECT 0.4 0.505 0.49 0.97 ;
  END
END SDFFX2H7R

MACRO SDFFX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFX3H7R 0 0 ;
  SIZE 8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 8 1.48 ;
        RECT 7.485 1.07 7.575 1.48 ;
        RECT 6.945 1.065 7.035 1.48 ;
        RECT 6.395 1.07 6.485 1.48 ;
        RECT 5.855 1.07 5.945 1.48 ;
        RECT 4.84 1.09 4.98 1.48 ;
        RECT 3.57 1.24 3.71 1.48 ;
        RECT 2.7 1.24 2.84 1.48 ;
        RECT 1.215 1.24 1.355 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 8 0.08 ;
        RECT 7.485 -0.08 7.575 0.345 ;
        RECT 6.945 -0.08 7.035 0.34 ;
        RECT 6.395 -0.08 6.485 0.345 ;
        RECT 5.855 -0.08 5.945 0.33 ;
        RECT 4.85 -0.08 4.99 0.275 ;
        RECT 3.575 -0.08 3.715 0.16 ;
        RECT 2.645 -0.08 2.785 0.16 ;
        RECT 1.025 -0.08 1.165 0.16 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 3.255 0.625 3.475 0.775 ;
      LAYER MET2 ;
        RECT 3.25 0.43 3.35 0.96 ;
      LAYER VIA1 ;
        RECT 3.255 0.655 3.345 0.745 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.26 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.655 0.21 6.745 1.145 ;
        RECT 6.125 0.805 6.745 0.895 ;
        RECT 6.215 0.435 6.745 0.525 ;
        RECT 6.215 0.225 6.305 0.525 ;
        RECT 6.125 0.805 6.215 1.13 ;
        RECT 6.1 0.225 6.305 0.315 ;
      LAYER MET2 ;
        RECT 6.65 0.425 6.75 0.96 ;
      LAYER VIA1 ;
        RECT 6.655 0.655 6.745 0.745 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.755 0.2 7.845 1.145 ;
        RECT 7.215 0.655 7.845 0.745 ;
        RECT 7.215 0.2 7.305 1.145 ;
      LAYER MET2 ;
        RECT 7.25 0.425 7.35 0.96 ;
      LAYER VIA1 ;
        RECT 7.255 0.655 7.345 0.745 ;
    END
  END QN
  PIN SE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.345 0.455 1.485 0.6 ;
        RECT 0.63 0.455 1.485 0.545 ;
        RECT 0.63 0.455 0.72 0.625 ;
      LAYER MET2 ;
        RECT 0.85 0.225 0.95 0.76 ;
      LAYER VIA1 ;
        RECT 0.855 0.455 0.945 0.545 ;
    END
  END SE
  PIN SI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.025 0.65 1.225 0.785 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END SI
  OBS
    LAYER MET1 ;
      RECT 5.495 0.55 5.585 1.005 ;
      RECT 6.025 0.625 6.34 0.715 ;
      RECT 4.885 0.55 5.675 0.64 ;
      RECT 5.585 0.295 5.675 0.64 ;
      RECT 6.025 0.455 6.115 0.715 ;
      RECT 5.585 0.455 6.115 0.545 ;
      RECT 5.07 1.14 5.765 1.23 ;
      RECT 5.675 0.8 5.765 1.23 ;
      RECT 5.07 0.91 5.16 1.23 ;
      RECT 4.1 0.91 5.16 1 ;
      RECT 4.1 0.35 4.19 1 ;
      RECT 5.675 0.8 5.935 0.89 ;
      RECT 5.845 0.655 5.935 0.89 ;
      RECT 4.1 0.35 4.245 0.44 ;
      RECT 5.25 0.73 5.34 1.005 ;
      RECT 4.36 0.73 5.34 0.82 ;
      RECT 4.36 0.17 4.45 0.82 ;
      RECT 2.305 0.25 2.395 0.575 ;
      RECT 4.36 0.365 5.43 0.455 ;
      RECT 5.34 0.295 5.43 0.455 ;
      RECT 3.496 0.25 3.915 0.34 ;
      RECT 2.305 0.25 2.97 0.34 ;
      RECT 3.454 0.191 3.496 0.319 ;
      RECT 3.416 0.25 3.915 0.279 ;
      RECT 3.825 0.17 4.45 0.26 ;
      RECT 2.88 0.231 3.534 0.26 ;
      RECT 2.88 0.17 3.454 0.26 ;
      RECT 3.89 1.14 4.325 1.23 ;
      RECT 1.945 1.125 2.51 1.215 ;
      RECT 2.42 1.06 3.98 1.15 ;
      RECT 1.945 0.48 2.035 1.215 ;
      RECT 3.89 0.43 3.98 1.23 ;
      RECT 3.29 0.43 3.98 0.52 ;
      RECT 3.29 0.355 3.38 0.52 ;
      RECT 3.06 0.88 3.765 0.97 ;
      RECT 3.675 0.64 3.765 0.97 ;
      RECT 3.06 0.35 3.15 0.97 ;
      RECT 2.545 0.475 3.15 0.565 ;
      RECT 2.125 0.85 2.92 0.94 ;
      RECT 2.83 0.665 2.92 0.94 ;
      RECT 2.125 0.24 2.215 0.94 ;
      RECT 2.83 0.665 2.97 0.755 ;
      RECT 0.705 1.06 1.855 1.15 ;
      RECT 1.765 0.17 1.855 1.15 ;
      RECT 1.765 0.17 1.91 0.345 ;
      RECT 0.505 0.25 1.35 0.34 ;
      RECT 1.26 0.17 1.91 0.26 ;
      RECT 0.4 0.88 1.665 0.97 ;
      RECT 1.575 0.35 1.665 0.97 ;
      RECT 0.84 0.75 0.93 0.97 ;
      RECT 0.4 0.505 0.49 0.97 ;
  END
END SDFFX3H7R

MACRO TBUFX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX0P5H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.04 0.935 1.13 1.48 ;
        RECT 0.32 0.945 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.04 -0.08 1.13 0.34 ;
        RECT 0.32 -0.08 0.41 0.335 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.625 0.37 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.905 0.45 1.175 0.55 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.66 0.935 0.925 1.025 ;
        RECT 0.625 0.235 0.925 0.35 ;
        RECT 0.66 0.235 0.75 1.025 ;
      LAYER MET2 ;
        RECT 0.65 0.18 0.75 0.56 ;
      LAYER VIA1 ;
        RECT 0.655 0.255 0.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.29 0.2 1.38 1.035 ;
      RECT 0.84 0.695 1.38 0.785 ;
      RECT 0.07 0.21 0.16 1.035 ;
      RECT 0.48 0.445 0.57 0.61 ;
      RECT 0.07 0.445 0.57 0.535 ;
  END
END TBUFX0P5H7R

MACRO TBUFX0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX0P7H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.04 0.935 1.13 1.48 ;
        RECT 0.32 0.945 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.04 -0.08 1.13 0.34 ;
        RECT 0.32 -0.08 0.41 0.335 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.625 0.37 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.905 0.45 1.175 0.55 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.66 0.935 0.925 1.025 ;
        RECT 0.625 0.255 0.925 0.345 ;
        RECT 0.66 0.255 0.75 1.025 ;
      LAYER MET2 ;
        RECT 0.65 0.18 0.75 0.56 ;
      LAYER VIA1 ;
        RECT 0.655 0.255 0.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.29 0.2 1.38 1.035 ;
      RECT 0.84 0.695 1.38 0.785 ;
      RECT 0.07 0.21 0.16 1.035 ;
      RECT 0.48 0.445 0.57 0.585 ;
      RECT 0.07 0.445 0.57 0.535 ;
  END
END TBUFX0P7H7R

MACRO TBUFX12H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX12H7R 0 0 ;
  SIZE 7 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7 1.48 ;
        RECT 6.775 1.035 6.865 1.48 ;
        RECT 6.235 1.15 6.375 1.48 ;
        RECT 5.705 1.15 5.845 1.48 ;
        RECT 5.175 1.15 5.315 1.48 ;
        RECT 4.62 1.035 4.71 1.48 ;
        RECT 2.855 1.095 2.995 1.48 ;
        RECT 2.355 1.095 2.495 1.48 ;
        RECT 1.855 1.095 1.995 1.48 ;
        RECT 1.34 1.195 1.48 1.48 ;
        RECT 0.85 1.05 0.94 1.48 ;
        RECT 0.32 1.05 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7 0.08 ;
        RECT 6.73 -0.08 6.82 0.365 ;
        RECT 6.175 -0.08 6.315 0.19 ;
        RECT 5.645 -0.08 5.785 0.19 ;
        RECT 5.11 -0.08 5.25 0.19 ;
        RECT 4.62 -0.08 4.71 0.35 ;
        RECT 4.08 -0.08 4.22 0.175 ;
        RECT 3.55 -0.08 3.69 0.175 ;
        RECT 3.015 -0.08 3.155 0.175 ;
        RECT 1.34 -0.08 1.48 0.175 ;
        RECT 0.85 -0.08 0.94 0.35 ;
        RECT 0.31 -0.08 0.45 0.185 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.005 0.655 1.345 0.745 ;
      LAYER MET2 ;
        RECT 1.05 0.425 1.15 0.96 ;
      LAYER VIA1 ;
        RECT 1.055 0.655 1.145 0.745 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.511 0.555 2.35 0.645 ;
        RECT 0.695 0.536 1.549 0.565 ;
        RECT 0.695 0.496 1.511 0.565 ;
        RECT 1.469 0.555 2.35 0.624 ;
        RECT 0.695 0.475 1.469 0.565 ;
        RECT 1.431 0.555 2.35 0.584 ;
        RECT 0.365 0.655 0.785 0.745 ;
        RECT 0.695 0.475 0.785 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.91 0.97 6.615 1.06 ;
        RECT 6.525 0.28 6.615 1.06 ;
        RECT 6.455 0.825 6.615 1.06 ;
        RECT 4.845 0.28 6.615 0.37 ;
      LAYER MET2 ;
        RECT 6.45 0.625 6.55 1.16 ;
      LAYER VIA1 ;
        RECT 6.455 0.855 6.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 3.604 0.96 4.314 1.05 ;
      RECT 4.224 0.265 4.314 1.05 ;
      RECT 4.224 0.51 6.315 0.6 ;
      RECT 2.825 0.265 4.485 0.355 ;
      RECT 1.075 0.265 1.75 0.355 ;
      RECT 1.66 0.17 1.75 0.355 ;
      RECT 2.814 0.221 2.825 0.35 ;
      RECT 2.768 0.193 2.814 0.321 ;
      RECT 2.73 0.246 2.863 0.279 ;
      RECT 1.66 0.17 2.768 0.26 ;
      RECT 3.13 1.14 4.494 1.23 ;
      RECT 4.404 0.74 4.494 1.23 ;
      RECT 3.13 0.915 3.22 1.23 ;
      RECT 1.075 1.015 1.72 1.105 ;
      RECT 1.63 0.915 1.72 1.105 ;
      RECT 1.63 0.915 3.51 1.005 ;
      RECT 3.42 0.445 3.51 1.005 ;
      RECT 4.404 0.74 6.245 0.83 ;
      RECT 2.673 0.445 3.51 0.535 ;
      RECT 2.662 0.401 2.673 0.53 ;
      RECT 2.616 0.373 2.662 0.501 ;
      RECT 2.578 0.426 2.711 0.459 ;
      RECT 1.885 0.35 2.616 0.44 ;
      RECT 0.07 0.275 0.16 1.095 ;
      RECT 0.6 0.835 0.69 1.08 ;
      RECT 0.07 0.835 1.444 0.925 ;
      RECT 0.07 0.835 1.49 0.902 ;
      RECT 1.406 0.816 1.544 0.844 ;
      RECT 1.49 0.743 1.506 0.871 ;
      RECT 3.24 0.64 3.33 0.825 ;
      RECT 1.444 0.774 3.33 0.825 ;
      RECT 1.506 0.735 3.33 0.825 ;
      RECT 0.07 0.275 0.715 0.365 ;
  END
END TBUFX12H7R

MACRO TBUFX16H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX16H7R 0 0 ;
  SIZE 9.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 9.8 1.48 ;
        RECT 9.281 1.055 9.371 1.48 ;
        RECT 8.756 1.095 8.896 1.48 ;
        RECT 8.256 1.095 8.396 1.48 ;
        RECT 7.746 1.095 7.886 1.48 ;
        RECT 7.246 1.095 7.386 1.48 ;
        RECT 6.771 1.055 6.861 1.48 ;
        RECT 4.155 1.075 4.295 1.48 ;
        RECT 3.655 1.075 3.795 1.48 ;
        RECT 3.155 1.075 3.295 1.48 ;
        RECT 2.655 1.075 2.795 1.48 ;
        RECT 2.14 1.205 2.28 1.48 ;
        RECT 1.61 1.205 1.75 1.48 ;
        RECT 1.12 1.05 1.21 1.48 ;
        RECT 0.57 1.05 0.66 1.48 ;
        RECT 0.07 1.035 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 9.8 0.08 ;
        RECT 9.29 -0.08 9.43 0.185 ;
        RECT 8.695 -0.08 8.835 0.185 ;
        RECT 8.135 -0.08 8.275 0.185 ;
        RECT 7.575 -0.08 7.715 0.185 ;
        RECT 7.015 -0.08 7.155 0.185 ;
        RECT 6.495 -0.08 6.585 0.35 ;
        RECT 5.94 -0.08 6.08 0.175 ;
        RECT 5.41 -0.08 5.55 0.175 ;
        RECT 4.88 -0.08 5.02 0.175 ;
        RECT 4.35 -0.08 4.49 0.175 ;
        RECT 2.14 -0.08 2.28 0.205 ;
        RECT 1.61 -0.08 1.75 0.205 ;
        RECT 1.12 -0.08 1.21 0.35 ;
        RECT 0.56 -0.08 0.7 0.225 ;
        RECT 0.07 -0.08 0.16 0.365 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.275 0.655 2.015 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.331 0.53 3.375 0.62 ;
        RECT 1.055 0.511 2.369 0.565 ;
        RECT 1.055 0.483 2.331 0.565 ;
        RECT 2.314 0.53 3.375 0.612 ;
        RECT 1.055 0.475 2.314 0.565 ;
        RECT 2.276 0.53 3.375 0.584 ;
        RECT 0.515 0.655 1.145 0.745 ;
        RECT 1.055 0.475 1.145 0.745 ;
      LAYER MET2 ;
        RECT 0.65 0.425 0.75 0.96 ;
      LAYER VIA1 ;
        RECT 0.655 0.655 0.745 0.745 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.735 0.275 9.71 0.365 ;
        RECT 7.021 0.915 9.146 1.005 ;
        RECT 9.055 0.275 9.146 1.005 ;
        RECT 8.031 0.915 8.121 1.08 ;
        RECT 7.521 0.915 7.611 1.06 ;
        RECT 7.021 0.915 7.111 1.08 ;
      LAYER MET2 ;
        RECT 9.05 0.225 9.15 0.76 ;
      LAYER VIA1 ;
        RECT 9.055 0.455 9.145 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 5.31 0.85 6.35 0.94 ;
      RECT 6.26 0.265 6.35 0.94 ;
      RECT 6.26 0.505 8.961 0.595 ;
      RECT 1.345 0.295 2.53 0.385 ;
      RECT 2.44 0.17 2.53 0.385 ;
      RECT 4.081 0.265 6.35 0.355 ;
      RECT 4.07 0.221 4.081 0.35 ;
      RECT 4.024 0.193 4.07 0.321 ;
      RECT 3.986 0.246 4.119 0.279 ;
      RECT 2.44 0.17 4.024 0.26 ;
      RECT 1.37 1.015 1.46 1.175 ;
      RECT 4.42 1.055 6.56 1.145 ;
      RECT 6.47 0.735 6.56 1.145 ;
      RECT 1.37 1.015 2.52 1.105 ;
      RECT 2.43 0.895 2.52 1.105 ;
      RECT 5.095 0.445 5.185 1.145 ;
      RECT 4.42 0.855 4.96 1.145 ;
      RECT 2.43 0.895 4.96 0.985 ;
      RECT 6.47 0.735 8.131 0.825 ;
      RECT 4.001 0.445 5.185 0.535 ;
      RECT 3.99 0.401 4.001 0.53 ;
      RECT 3.944 0.373 3.99 0.501 ;
      RECT 3.906 0.426 4.039 0.459 ;
      RECT 2.665 0.35 3.944 0.44 ;
      RECT 0.85 0.835 0.94 1.025 ;
      RECT 0.32 0.315 0.41 1.025 ;
      RECT 0.32 0.835 2.204 0.925 ;
      RECT 0.32 0.835 2.25 0.902 ;
      RECT 2.166 0.816 2.291 0.859 ;
      RECT 2.204 0.774 2.329 0.819 ;
      RECT 2.25 0.73 2.291 0.859 ;
      RECT 2.291 0.71 4.34 0.8 ;
      RECT 4.25 0.625 5.005 0.715 ;
      RECT 0.32 0.315 0.965 0.405 ;
  END
END TBUFX16H7R

MACRO TBUFX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX1H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.04 0.895 1.13 1.48 ;
        RECT 0.305 0.91 0.445 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.04 -0.08 1.13 0.335 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.625 0.39 0.82 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.9 0.455 1.2 0.545 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.66 0.895 0.925 0.985 ;
        RECT 0.625 0.255 0.925 0.345 ;
        RECT 0.66 0.255 0.75 0.985 ;
      LAYER MET2 ;
        RECT 0.65 0.18 0.75 0.56 ;
      LAYER VIA1 ;
        RECT 0.655 0.255 0.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.29 0.195 1.38 0.995 ;
      RECT 0.84 0.685 1.38 0.775 ;
      RECT 0.07 0.205 0.16 0.995 ;
      RECT 0.48 0.445 0.57 0.645 ;
      RECT 0.07 0.445 0.57 0.535 ;
  END
END TBUFX1H7R

MACRO TBUFX1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX1P4H7R 0 0 ;
  SIZE 1.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.6 1.48 ;
        RECT 1.04 0.895 1.13 1.48 ;
        RECT 0.35 1.029 0.44 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.6 0.08 ;
        RECT 1.04 -0.08 1.13 0.335 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.62 0.385 0.82 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.9 0.455 1.2 0.545 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.66 0.915 0.925 1.005 ;
        RECT 0.625 0.255 0.925 0.345 ;
        RECT 0.66 0.255 0.75 1.005 ;
      LAYER MET2 ;
        RECT 0.65 0.18 0.75 0.56 ;
      LAYER VIA1 ;
        RECT 0.655 0.255 0.745 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.29 0.195 1.38 0.995 ;
      RECT 0.855 0.685 1.38 0.775 ;
      RECT 0.07 0.205 0.16 0.99 ;
      RECT 0.48 0.44 0.57 0.65 ;
      RECT 0.07 0.44 0.57 0.53 ;
  END
END TBUFX1P4H7R

MACRO TBUFX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX2H7R 0 0 ;
  SIZE 2.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.2 1.48 ;
        RECT 1.755 0.95 1.895 1.48 ;
        RECT 0.79 1.09 0.93 1.48 ;
        RECT 0.32 0.93 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.2 0.08 ;
        RECT 1.755 -0.08 1.895 0.335 ;
        RECT 0.79 -0.08 0.93 0.295 ;
        RECT 0.295 -0.08 0.435 0.335 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.4 0.605 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.795 0.425 1.945 0.605 ;
      LAYER MET2 ;
        RECT 1.85 0.225 1.95 0.76 ;
      LAYER VIA1 ;
        RECT 1.855 0.455 1.945 0.545 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.255 0.35 1.405 0.985 ;
      LAYER MET2 ;
        RECT 1.25 0.23 1.35 0.76 ;
      LAYER VIA1 ;
        RECT 1.255 0.455 1.345 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.035 0.22 2.125 1.025 ;
      RECT 1.495 0.7 2.125 0.84 ;
      RECT 1.05 1.115 1.655 1.205 ;
      RECT 1.515 0.95 1.655 1.205 ;
      RECT 1.05 0.91 1.14 1.205 ;
      RECT 0.525 0.91 1.14 1 ;
      RECT 0.55 0.385 1.135 0.475 ;
      RECT 1.045 0.17 1.135 0.475 ;
      RECT 1.54 0.17 1.63 0.45 ;
      RECT 0.55 0.31 0.64 0.475 ;
      RECT 1.045 0.17 1.63 0.26 ;
      RECT 0.07 0.22 0.16 1.03 ;
      RECT 0.07 0.71 0.915 0.8 ;
  END
END TBUFX2H7R

MACRO TBUFX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX3H7R 0 0 ;
  SIZE 3 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3 1.48 ;
        RECT 2.55 1.05 2.64 1.48 ;
        RECT 1.025 1.105 1.115 1.48 ;
        RECT 0.345 1.12 0.485 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3 0.08 ;
        RECT 2.55 -0.08 2.64 0.33 ;
        RECT 1.545 -0.08 1.685 0.175 ;
        RECT 0.355 -0.08 0.495 0.335 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.44 0.625 0.575 0.825 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.772 0.555 0.99 0.645 ;
        RECT 0.68 0.536 0.81 0.576 ;
        RECT 0.68 0.494 0.772 0.576 ;
        RECT 0.726 0.555 0.99 0.622 ;
        RECT 0.255 0.448 0.726 0.515 ;
        RECT 0.255 0.425 0.68 0.515 ;
        RECT 0.642 0.494 0.772 0.534 ;
        RECT 0.255 0.425 0.345 0.645 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.8 0.28 2.89 1.04 ;
        RECT 2.3 0.87 2.89 0.96 ;
        RECT 2.3 0.455 2.89 0.545 ;
        RECT 2.3 0.87 2.39 1.04 ;
        RECT 2.3 0.28 2.39 0.545 ;
      LAYER MET2 ;
        RECT 2.65 0.23 2.75 0.76 ;
      LAYER VIA1 ;
        RECT 2.655 0.455 2.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.33 1.14 2.21 1.23 ;
      RECT 2.12 0.265 2.21 1.23 ;
      RECT 0.635 1.12 0.777 1.21 ;
      RECT 0.635 1.12 0.823 1.187 ;
      RECT 1.33 0.925 1.42 1.23 ;
      RECT 0.739 1.101 0.869 1.141 ;
      RECT 0.777 1.059 0.869 1.141 ;
      RECT 0.777 1.059 0.915 1.095 ;
      RECT 0.823 1.013 0.934 1.063 ;
      RECT 0.823 1.013 0.972 1.034 ;
      RECT 0.934 0.925 1.42 1.015 ;
      RECT 0.869 0.967 1.42 1.015 ;
      RECT 0.915 0.934 0.934 1.063 ;
      RECT 1.465 0.265 2.21 0.355 ;
      RECT 1.433 0.211 1.465 0.339 ;
      RECT 1.395 0.265 2.21 0.304 ;
      RECT 0.935 0.195 1.433 0.285 ;
      RECT 0.935 0.246 1.503 0.285 ;
      RECT 1.53 0.945 2.03 1.035 ;
      RECT 1.94 0.445 2.03 1.035 ;
      RECT 1.386 0.445 2.03 0.535 ;
      RECT 1.354 0.391 1.386 0.519 ;
      RECT 1.316 0.445 2.03 0.484 ;
      RECT 0.855 0.375 1.354 0.465 ;
      RECT 0.855 0.426 1.424 0.465 ;
      RECT 0.809 0.314 0.855 0.442 ;
      RECT 0.763 0.268 0.809 0.396 ;
      RECT 0.763 0.356 0.893 0.396 ;
      RECT 0.725 0.314 0.855 0.354 ;
      RECT 0.615 0.245 0.763 0.335 ;
      RECT 0.07 0.94 0.662 1.03 ;
      RECT 0.07 0.94 0.708 1.007 ;
      RECT 0.624 0.921 0.754 0.961 ;
      RECT 0.07 0.295 0.16 1.03 ;
      RECT 0.662 0.879 0.754 0.961 ;
      RECT 0.708 0.833 0.8 0.915 ;
      RECT 0.754 0.787 0.867 0.844 ;
      RECT 0.8 0.749 0.829 0.878 ;
      RECT 0.829 0.735 1.77 0.825 ;
  END
END TBUFX3H7R

MACRO TBUFX4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX4H7R 0 0 ;
  SIZE 3.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.4 1.48 ;
        RECT 2.964 1.05 3.054 1.48 ;
        RECT 0.985 1.09 1.125 1.48 ;
        RECT 0.295 1.09 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.4 0.08 ;
        RECT 2.972 -0.08 3.062 0.33 ;
        RECT 2.472 -0.08 2.562 0.33 ;
        RECT 2.202 -0.08 2.342 0.195 ;
        RECT 1.576 -0.08 1.721 0.16 ;
        RECT 0.32 -0.08 0.41 0.335 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 0.625 0.6 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.727 0.53 1.17 0.62 ;
        RECT 0.622 0.511 0.765 0.534 ;
        RECT 0.255 0.481 0.727 0.515 ;
        RECT 0.706 0.53 1.17 0.61 ;
        RECT 0.255 0.448 0.706 0.515 ;
        RECT 0.66 0.53 1.17 0.576 ;
        RECT 0.255 0.425 0.66 0.515 ;
        RECT 0.255 0.425 0.345 0.68 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.214 0.225 3.345 1.15 ;
        RECT 2.714 0.87 3.345 0.96 ;
        RECT 2.722 0.42 3.345 0.51 ;
        RECT 2.722 0.27 2.812 0.51 ;
        RECT 2.714 0.87 2.804 1.015 ;
      LAYER MET2 ;
        RECT 3.25 0.18 3.35 0.56 ;
      LAYER VIA1 ;
        RECT 3.255 0.255 3.345 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.285 1.14 2.624 1.23 ;
      RECT 2.534 0.593 2.624 1.23 ;
      RECT 0.555 1.09 0.764 1.18 ;
      RECT 0.555 1.09 0.81 1.157 ;
      RECT 1.285 0.9 1.375 1.23 ;
      RECT 0.726 1.071 0.856 1.111 ;
      RECT 0.764 1.029 0.856 1.111 ;
      RECT 0.764 1.029 0.902 1.065 ;
      RECT 0.81 0.983 0.916 1.035 ;
      RECT 0.81 0.983 0.954 1.009 ;
      RECT 0.916 0.9 1.375 0.99 ;
      RECT 0.856 0.937 1.375 0.99 ;
      RECT 0.902 0.907 0.916 1.035 ;
      RECT 2.524 0.52 2.534 0.648 ;
      RECT 2.478 0.492 2.524 0.62 ;
      RECT 2.478 0.548 2.58 0.62 ;
      RECT 2.432 0.446 2.478 0.574 ;
      RECT 2.386 0.4 2.432 0.528 ;
      RECT 2.34 0.354 2.386 0.482 ;
      RECT 2.294 0.308 2.34 0.436 ;
      RECT 2.256 0.354 2.386 0.394 ;
      RECT 1.531 0.285 2.294 0.375 ;
      RECT 1.5 0.231 1.531 0.36 ;
      RECT 1.454 0.193 1.5 0.321 ;
      RECT 1.454 0.266 1.569 0.321 ;
      RECT 1.416 0.17 1.454 0.279 ;
      RECT 0.915 0.17 1.454 0.26 ;
      RECT 1.588 0.95 2.405 1.04 ;
      RECT 1.972 0.465 2.062 1.04 ;
      RECT 1.972 0.67 2.419 0.76 ;
      RECT 1.26 0.465 2.062 0.555 ;
      RECT 1.26 0.35 1.375 0.555 ;
      RECT 0.83 0.35 1.375 0.44 ;
      RECT 0.794 0.294 0.83 0.422 ;
      RECT 0.748 0.253 0.794 0.381 ;
      RECT 0.748 0.331 0.868 0.381 ;
      RECT 0.71 0.23 0.748 0.339 ;
      RECT 0.6 0.23 0.748 0.32 ;
      RECT 0.07 0.31 0.16 1.03 ;
      RECT 0.07 0.91 0.677 1 ;
      RECT 0.07 0.91 0.723 0.977 ;
      RECT 0.639 0.891 0.769 0.931 ;
      RECT 0.677 0.849 0.769 0.931 ;
      RECT 0.677 0.849 0.815 0.885 ;
      RECT 0.723 0.803 0.839 0.85 ;
      RECT 1.64 0.685 1.73 0.825 ;
      RECT 1.44 0.685 1.53 0.825 ;
      RECT 0.769 0.757 0.877 0.819 ;
      RECT 0.815 0.722 0.839 0.85 ;
      RECT 0.839 0.71 1.755 0.8 ;
  END
END TBUFX4H7R

MACRO TBUFX6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX6H7R 0 0 ;
  SIZE 5.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.2 1.48 ;
        RECT 4.988 1.045 5.078 1.48 ;
        RECT 4.488 1.06 4.578 1.48 ;
        RECT 3.988 1.045 4.078 1.48 ;
        RECT 2.275 1.12 2.365 1.48 ;
        RECT 1.73 1.125 1.82 1.48 ;
        RECT 1.12 1.196 1.26 1.48 ;
        RECT 0.32 1.053 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.2 0.08 ;
        RECT 4.92 -0.08 5.01 0.375 ;
        RECT 4.42 -0.08 4.51 0.36 ;
        RECT 3.92 -0.08 4.01 0.375 ;
        RECT 3.175 -0.08 3.315 0.16 ;
        RECT 2.555 -0.08 2.695 0.16 ;
        RECT 1.135 -0.08 1.275 0.17 ;
        RECT 0.34 -0.08 0.48 0.175 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.035 0.655 1.375 0.745 ;
      LAYER MET2 ;
        RECT 1.25 0.43 1.35 0.96 ;
      LAYER VIA1 ;
        RECT 1.255 0.655 1.345 0.745 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.52 0.58 2.16 0.67 ;
        RECT 1.41 0.568 1.59 0.583 ;
        RECT 1.41 0.533 1.566 0.583 ;
        RECT 0.25 0.505 1.52 0.56 ;
        RECT 1.511 0.58 2.16 0.666 ;
        RECT 0.25 0.478 1.511 0.56 ;
        RECT 1.465 0.58 2.16 0.638 ;
        RECT 0.25 0.455 1.465 0.56 ;
        RECT 1.456 0.58 2.16 0.611 ;
      LAYER MET2 ;
        RECT 0.45 0.23 0.55 0.76 ;
      LAYER VIA1 ;
        RECT 0.455 0.455 0.545 0.545 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.738 0.325 4.828 1.037 ;
        RECT 4.238 0.88 4.828 0.97 ;
        RECT 4.17 0.455 4.828 0.545 ;
        RECT 4.67 0.325 4.828 0.545 ;
        RECT 4.238 0.88 4.328 1.035 ;
        RECT 4.17 0.325 4.26 0.545 ;
      LAYER MET2 ;
        RECT 4.65 0.225 4.75 0.76 ;
      LAYER VIA1 ;
        RECT 4.655 0.455 4.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.95 1.14 3.83 1.23 ;
      RECT 3.74 0.28 3.83 1.23 ;
      RECT 3.45 0.94 3.54 1.23 ;
      RECT 2.95 0.94 3.04 1.23 ;
      RECT 0.855 1.016 1.621 1.106 ;
      RECT 0.855 1.016 1.697 1.049 ;
      RECT 1.659 0.94 3.04 1.03 ;
      RECT 1.583 0.997 3.04 1.03 ;
      RECT 1.621 0.959 1.659 1.087 ;
      RECT 3.74 0.805 3.933 0.895 ;
      RECT 2.478 0.25 3.829 0.34 ;
      RECT 2.436 0.191 2.478 0.319 ;
      RECT 2.398 0.25 3.829 0.279 ;
      RECT 1.675 0.17 2.436 0.26 ;
      RECT 1.675 0.231 2.516 0.26 ;
      RECT 3.2 0.43 3.29 1.045 ;
      RECT 3.56 0.43 3.65 0.746 ;
      RECT 2.395 0.43 3.65 0.52 ;
      RECT 2.353 0.371 2.395 0.499 ;
      RECT 2.315 0.43 3.65 0.459 ;
      RECT 1.592 0.35 2.353 0.44 ;
      RECT 1.592 0.411 2.433 0.44 ;
      RECT 1.555 0.293 1.592 0.422 ;
      RECT 1.517 0.275 1.555 0.384 ;
      RECT 0.855 0.275 1.555 0.365 ;
      RECT 0.855 0.331 1.63 0.365 ;
      RECT 0.63 0.835 0.72 1.155 ;
      RECT 0.07 0.275 0.16 1.155 ;
      RECT 0.07 0.835 1.537 0.925 ;
      RECT 0.07 0.835 1.574 0.907 ;
      RECT 0.07 0.835 1.612 0.869 ;
      RECT 2.513 0.66 2.603 0.85 ;
      RECT 1.499 0.816 2.603 0.85 ;
      RECT 1.574 0.76 2.603 0.85 ;
      RECT 1.537 0.778 2.603 0.85 ;
      RECT 2.513 0.66 3.11 0.75 ;
      RECT 0.07 0.275 0.745 0.365 ;
  END
END TBUFX6H7R

MACRO TBUFX8H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX8H7R 0 0 ;
  SIZE 5.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.2 1.48 ;
        RECT 4.712 1.095 4.852 1.48 ;
        RECT 4.212 1.095 4.352 1.48 ;
        RECT 3.737 1.055 3.827 1.48 ;
        RECT 2.185 1.195 2.325 1.48 ;
        RECT 1.655 1.195 1.795 1.48 ;
        RECT 1.125 1.195 1.265 1.48 ;
        RECT 0.56 1.075 0.7 1.48 ;
        RECT 0.06 1.075 0.2 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.2 0.08 ;
        RECT 4.7 -0.08 4.84 0.305 ;
        RECT 4.2 -0.08 4.34 0.305 ;
        RECT 3.725 -0.08 3.815 0.33 ;
        RECT 3.19 -0.08 3.33 0.175 ;
        RECT 2.66 -0.08 2.8 0.175 ;
        RECT 1.14 -0.08 1.28 0.16 ;
        RECT 0.585 -0.08 0.675 0.335 ;
        RECT 0.085 -0.08 0.175 0.35 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.745 0.655 1.045 0.745 ;
      LAYER MET2 ;
        RECT 0.85 0.425 0.95 0.96 ;
      LAYER VIA1 ;
        RECT 0.855 0.655 0.945 0.745 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.319 0.625 2.12 0.715 ;
        RECT 1.207 0.606 1.357 0.626 ;
        RECT 1.207 0.577 1.319 0.626 ;
        RECT 1.299 0.625 2.12 0.705 ;
        RECT 1.169 0.544 1.299 0.584 ;
        RECT 1.253 0.625 2.12 0.672 ;
        RECT 0.515 0.498 1.253 0.565 ;
        RECT 0.515 0.475 1.207 0.565 ;
        RECT 0.38 0.655 0.605 0.745 ;
        RECT 0.515 0.475 0.605 0.745 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.962 0.911 5.102 1.001 ;
        RECT 5.012 0.295 5.102 1.001 ;
        RECT 3.975 0.455 5.102 0.545 ;
        RECT 4.975 0.295 5.102 0.545 ;
        RECT 4.475 0.31 4.565 0.545 ;
        RECT 3.975 0.31 4.065 0.545 ;
      LAYER MET2 ;
        RECT 4.9 0.225 5 0.76 ;
      LAYER VIA1 ;
        RECT 4.905 0.455 4.995 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 3.17 0.355 3.26 1 ;
      RECT 3.505 0.525 3.781 0.615 ;
      RECT 3.505 0.355 3.595 0.615 ;
      RECT 2.403 0.355 3.595 0.445 ;
      RECT 2.367 0.299 2.403 0.427 ;
      RECT 2.321 0.258 2.367 0.386 ;
      RECT 2.321 0.336 2.441 0.386 ;
      RECT 2.283 0.235 2.321 0.344 ;
      RECT 0.81 0.25 1.356 0.34 ;
      RECT 0.81 0.25 1.371 0.333 ;
      RECT 1.333 0.235 2.321 0.325 ;
      RECT 1.318 0.242 2.321 0.325 ;
      RECT 2.99 1.09 3.51 1.18 ;
      RECT 3.42 0.766 3.51 1.18 ;
      RECT 0.81 1.015 3.08 1.105 ;
      RECT 2.99 0.535 3.08 1.18 ;
      RECT 3.42 0.766 3.705 0.856 ;
      RECT 2.252 0.535 3.08 0.625 ;
      RECT 2.236 0.469 2.252 0.617 ;
      RECT 2.19 0.438 2.236 0.586 ;
      RECT 2.178 0.529 2.31 0.557 ;
      RECT 2.178 0.5 2.298 0.557 ;
      RECT 2.132 0.5 2.298 0.528 ;
      RECT 1.68 0.415 2.19 0.505 ;
      RECT 0.2 0.885 0.658 0.975 ;
      RECT 0.2 0.885 0.67 0.969 ;
      RECT 0.2 0.885 0.708 0.944 ;
      RECT 0.2 0.885 2.361 0.925 ;
      RECT 0.62 0.866 2.407 0.902 ;
      RECT 0.2 0.455 0.29 0.975 ;
      RECT 0.658 0.841 2.407 0.902 ;
      RECT 0.67 0.835 2.443 0.861 ;
      RECT 2.323 0.816 2.443 0.861 ;
      RECT 2.361 0.774 2.481 0.824 ;
      RECT 2.407 0.733 2.443 0.861 ;
      RECT 2.443 0.715 2.9 0.805 ;
      RECT 0.2 0.455 0.425 0.545 ;
      RECT 0.335 0.325 0.425 0.545 ;
  END
END TBUFX8H7R

MACRO TIEHIH7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TIEHIH7R 0 0 ;
  SIZE 0.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.8 1.48 ;
        RECT 0.575 1.055 0.665 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.8 0.08 ;
        RECT 0.57 -0.08 0.66 0.345 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 1.025 0.435 1.175 ;
      LAYER MET2 ;
        RECT 0.25 0.84 0.35 1.22 ;
      LAYER VIA1 ;
        RECT 0.255 1.055 0.345 1.145 ;
    END
  END Z
  OBS
    LAYER MET1 ;
      RECT 0.195 0.46 0.535 0.55 ;
      RECT 0.32 0.205 0.41 0.55 ;
  END
END TIEHIH7R

MACRO TIELOH7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TIELOH7R 0 0 ;
  SIZE 0.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 0.8 1.48 ;
        RECT 0.575 1.055 0.665 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 0.8 0.08 ;
        RECT 0.57 -0.08 0.66 0.345 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.22 0.41 0.395 ;
      LAYER MET2 ;
        RECT 0.25 0.18 0.35 0.56 ;
      LAYER VIA1 ;
        RECT 0.255 0.255 0.345 0.345 ;
    END
  END Z
  OBS
    LAYER MET1 ;
      RECT 0.32 0.73 0.41 1.155 ;
      RECT 0.195 0.73 0.535 0.82 ;
  END
END TIELOH7R

MACRO TINVX0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TINVX0P5H7R 0 0 ;
  SIZE 1.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.2 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.2 0.08 ;
        RECT 0.295 -0.08 0.435 0.325 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.825 0.545 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.42 0.805 0.545 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.805 1.06 1.145 1.15 ;
        RECT 1.055 0.235 1.145 1.15 ;
        RECT 0.815 0.235 1.145 0.325 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 1.035 0.16 1.175 ;
      RECT 0.045 0.21 0.135 1.175 ;
      RECT 0.69 0.635 0.78 0.945 ;
      RECT 0.045 0.635 0.78 0.725 ;
      RECT 0.045 0.21 0.16 0.35 ;
  END
END TINVX0P5H7R

MACRO TINVX0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TINVX0P7H7R 0 0 ;
  SIZE 1.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.2 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.2 0.08 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 0.635 0.6 0.77 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.455 0.82 0.545 ;
        RECT 0.225 0.455 0.315 0.595 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.795 1.04 1 1.13 ;
        RECT 0.91 0.245 1 1.13 ;
        RECT 0.795 0.245 1 0.345 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.56 ;
      LAYER VIA1 ;
        RECT 0.855 0.255 0.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.86 0.16 1.155 ;
      RECT 0.045 0.86 0.795 0.95 ;
      RECT 0.705 0.773 0.795 0.95 ;
      RECT 0.045 0.23 0.135 1.155 ;
      RECT 0.045 0.23 0.185 0.32 ;
  END
END TINVX0P7H7R

MACRO TINVX12H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TINVX12H7R 0 0 ;
  SIZE 9.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 9.8 1.48 ;
        RECT 9.25 1.07 9.34 1.48 ;
        RECT 8.74 1.07 8.83 1.48 ;
        RECT 8.15 1.225 8.29 1.48 ;
        RECT 7.61 1.055 7.7 1.48 ;
        RECT 5.445 1.07 5.585 1.48 ;
        RECT 4.97 1.07 5.06 1.48 ;
        RECT 4.47 1.07 4.56 1.48 ;
        RECT 3.97 1.07 4.06 1.48 ;
        RECT 3.25 1.07 3.34 1.48 ;
        RECT 2.75 1.07 2.84 1.48 ;
        RECT 2.25 1.07 2.34 1.48 ;
        RECT 1.635 0.87 1.725 1.48 ;
        RECT 1.07 0.87 1.16 1.48 ;
        RECT 0.57 0.87 0.66 1.48 ;
        RECT 0.07 0.855 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 9.8 0.08 ;
        RECT 9.63 -0.08 9.72 0.345 ;
        RECT 9.13 -0.08 9.22 0.33 ;
        RECT 8.63 -0.08 8.72 0.33 ;
        RECT 8.13 -0.08 8.22 0.33 ;
        RECT 7.63 -0.08 7.72 0.345 ;
        RECT 7.125 -0.08 7.265 0.305 ;
        RECT 6.625 -0.08 6.765 0.305 ;
        RECT 6.06 -0.08 6.2 0.175 ;
        RECT 4.04 -0.08 4.13 0.345 ;
        RECT 3.32 -0.08 3.41 0.33 ;
        RECT 2.82 -0.08 2.91 0.33 ;
        RECT 2.32 -0.08 2.41 0.33 ;
        RECT 1.82 -0.08 1.91 0.33 ;
        RECT 1.32 -0.08 1.41 0.33 ;
        RECT 0.82 -0.08 0.91 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.425 0.435 0.575 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.375 0.61 3.575 0.745 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 8.49 0.89 9.615 0.98 ;
        RECT 7.88 0.42 9.47 0.51 ;
        RECT 9.38 0.295 9.47 0.51 ;
        RECT 9.055 0.42 9.145 0.98 ;
        RECT 8.88 0.295 8.97 0.51 ;
        RECT 7.835 1.045 8.58 1.135 ;
        RECT 8.49 0.89 8.58 1.135 ;
        RECT 8.38 0.295 8.47 0.51 ;
        RECT 7.88 0.295 7.97 0.51 ;
      LAYER MET2 ;
        RECT 9.05 0.425 9.15 0.96 ;
      LAYER VIA1 ;
        RECT 9.055 0.655 9.145 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 4.72 0.865 4.81 1.195 ;
      RECT 2 0.855 2.09 1.195 ;
      RECT 5.7 0.865 5.79 1.18 ;
      RECT 5.22 0.865 5.31 1.18 ;
      RECT 4.22 0.865 4.31 1.18 ;
      RECT 3 0.855 3.09 1.17 ;
      RECT 2.5 0.855 2.59 1.17 ;
      RECT 3.43 1.075 3.88 1.165 ;
      RECT 3.79 0.961 3.88 1.165 ;
      RECT 3.43 0.855 3.52 1.165 ;
      RECT 3.836 0.916 3.947 0.974 ;
      RECT 3.88 0.879 3.909 1.008 ;
      RECT 7.765 0.71 7.855 0.955 ;
      RECT 2 0.855 3.52 0.945 ;
      RECT 3.909 0.865 7.855 0.955 ;
      RECT 6.117 0.445 6.207 0.955 ;
      RECT 7.765 0.71 8.905 0.8 ;
      RECT 4.52 0.445 6.207 0.535 ;
      RECT 5.52 0.36 5.61 0.535 ;
      RECT 5.02 0.36 5.11 0.535 ;
      RECT 4.52 0.36 4.61 0.535 ;
      RECT 7.4 0.59 7.635 0.68 ;
      RECT 7.4 0.35 7.49 0.68 ;
      RECT 3.86 0.435 4.36 0.525 ;
      RECT 4.27 0.17 4.36 0.525 ;
      RECT 2.07 0.42 3.59 0.51 ;
      RECT 3.5 0.19 3.59 0.51 ;
      RECT 6.4 0.395 7.49 0.485 ;
      RECT 3.86 0.19 3.95 0.525 ;
      RECT 3.07 0.37 3.16 0.51 ;
      RECT 2.57 0.37 2.66 0.51 ;
      RECT 2.07 0.37 2.16 0.51 ;
      RECT 6.4 0.265 6.49 0.485 ;
      RECT 5.77 0.265 6.49 0.355 ;
      RECT 5.27 0.17 5.36 0.33 ;
      RECT 4.77 0.17 4.86 0.33 ;
      RECT 3.5 0.19 3.95 0.28 ;
      RECT 5.77 0.17 5.86 0.355 ;
      RECT 4.27 0.17 5.86 0.26 ;
      RECT 3.61 0.822 3.7 0.985 ;
      RECT 3.61 0.822 3.746 0.86 ;
      RECT 3.68 0.37 3.77 0.825 ;
      RECT 3.656 0.787 3.77 0.825 ;
      RECT 3.68 0.625 6.004 0.715 ;
      RECT 1.32 0.665 1.41 1.15 ;
      RECT 0.82 0.665 0.91 1.15 ;
      RECT 0.32 0.665 0.41 1.15 ;
      RECT 0.07 0.665 1.66 0.755 ;
      RECT 1.57 0.37 1.66 0.755 ;
      RECT 1.57 0.625 3.255 0.715 ;
      RECT 1.07 0.37 1.16 0.755 ;
      RECT 0.57 0.27 0.66 0.755 ;
      RECT 0.07 0.255 0.16 0.755 ;
      RECT 9.57 0.525 9.72 0.705 ;
      RECT 5.925 1.08 7.495 1.17 ;
  END
END TINVX12H7R

MACRO TINVX16H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TINVX16H7R 0 0 ;
  SIZE 12.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 12.8 1.48 ;
        RECT 12.61 1.055 12.7 1.48 ;
        RECT 12.085 1.095 12.225 1.48 ;
        RECT 11.585 1.095 11.725 1.48 ;
        RECT 11.075 1.095 11.215 1.48 ;
        RECT 10.51 1.225 10.65 1.48 ;
        RECT 9.97 1.055 10.06 1.48 ;
        RECT 7.31 1.07 7.4 1.48 ;
        RECT 6.81 1.07 6.9 1.48 ;
        RECT 6.31 1.07 6.4 1.48 ;
        RECT 5.81 1.07 5.9 1.48 ;
        RECT 4.97 1.07 5.06 1.48 ;
        RECT 4.25 1.07 4.34 1.48 ;
        RECT 3.75 1.07 3.84 1.48 ;
        RECT 3.25 1.07 3.34 1.48 ;
        RECT 2.75 1.07 2.84 1.48 ;
        RECT 2.07 0.87 2.16 1.48 ;
        RECT 1.57 0.87 1.66 1.48 ;
        RECT 1.07 0.87 1.16 1.48 ;
        RECT 0.57 0.87 0.66 1.48 ;
        RECT 0.07 0.855 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 12.8 0.08 ;
        RECT 12.49 -0.08 12.58 0.345 ;
        RECT 11.99 -0.08 12.08 0.33 ;
        RECT 11.49 -0.08 11.58 0.33 ;
        RECT 10.99 -0.08 11.08 0.33 ;
        RECT 10.49 -0.08 10.58 0.33 ;
        RECT 9.99 -0.08 10.08 0.345 ;
        RECT 9.485 -0.08 9.625 0.305 ;
        RECT 8.985 -0.08 9.125 0.305 ;
        RECT 8.485 -0.08 8.625 0.305 ;
        RECT 7.92 -0.08 8.06 0.175 ;
        RECT 5.04 -0.08 5.13 0.33 ;
        RECT 4.32 -0.08 4.41 0.33 ;
        RECT 3.795 -0.08 3.935 0.305 ;
        RECT 3.295 -0.08 3.435 0.305 ;
        RECT 2.795 -0.08 2.935 0.305 ;
        RECT 2.32 -0.08 2.41 0.33 ;
        RECT 1.82 -0.08 1.91 0.33 ;
        RECT 1.32 -0.08 1.41 0.33 ;
        RECT 0.82 -0.08 0.91 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.255 0.425 0.435 0.575 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.255 0.625 4.52 0.775 ;
      LAYER MET2 ;
        RECT 4.25 0.425 4.35 0.96 ;
      LAYER VIA1 ;
        RECT 4.255 0.655 4.345 0.745 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 10.85 0.915 12.475 1.005 ;
        RECT 10.24 0.42 12.33 0.51 ;
        RECT 12.24 0.31 12.33 0.51 ;
        RECT 12.055 0.42 12.145 1.005 ;
        RECT 11.74 0.31 11.83 0.51 ;
        RECT 11.24 0.295 11.33 0.51 ;
        RECT 10.195 1.045 10.94 1.135 ;
        RECT 10.85 0.915 10.94 1.135 ;
        RECT 10.74 0.295 10.83 0.51 ;
        RECT 10.24 0.295 10.33 0.51 ;
      LAYER MET2 ;
        RECT 12.05 0.425 12.15 0.96 ;
      LAYER VIA1 ;
        RECT 12.055 0.655 12.145 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 5.15 1.105 5.65 1.195 ;
      RECT 5.56 0.855 5.65 1.195 ;
      RECT 4 0.88 4.09 1.195 ;
      RECT 3.5 0.88 3.59 1.195 ;
      RECT 3 0.88 3.09 1.195 ;
      RECT 2.5 0.855 2.59 1.195 ;
      RECT 7.56 0.86 7.65 1.175 ;
      RECT 7.06 0.86 7.15 1.175 ;
      RECT 6.56 0.86 6.65 1.175 ;
      RECT 6.06 0.86 6.15 1.175 ;
      RECT 4.43 1.04 4.88 1.13 ;
      RECT 4.79 0.89 4.88 1.13 ;
      RECT 5.15 0.89 5.24 1.195 ;
      RECT 4.43 0.88 4.52 1.13 ;
      RECT 4.79 0.89 5.24 0.98 ;
      RECT 2.5 0.88 4.52 0.97 ;
      RECT 5.56 0.86 10.255 0.95 ;
      RECT 10.165 0.72 10.255 0.95 ;
      RECT 7.977 0.445 8.067 0.95 ;
      RECT 10.165 0.72 11.815 0.81 ;
      RECT 5.88 0.445 8.067 0.535 ;
      RECT 7.38 0.36 7.47 0.535 ;
      RECT 6.88 0.36 6.97 0.535 ;
      RECT 6.38 0.36 6.47 0.535 ;
      RECT 5.88 0.36 5.97 0.535 ;
      RECT 9.76 0.59 9.955 0.68 ;
      RECT 9.76 0.355 9.85 0.68 ;
      RECT 4.86 0.42 5.31 0.51 ;
      RECT 5.22 0.17 5.31 0.51 ;
      RECT 4.14 0.42 4.59 0.51 ;
      RECT 4.5 0.19 4.59 0.51 ;
      RECT 8.26 0.395 9.85 0.485 ;
      RECT 2.545 0.395 4.23 0.485 ;
      RECT 4.86 0.19 4.95 0.51 ;
      RECT 8.26 0.265 8.35 0.485 ;
      RECT 7.63 0.265 8.35 0.355 ;
      RECT 5.63 0.17 5.72 0.345 ;
      RECT 7.13 0.17 7.22 0.33 ;
      RECT 6.63 0.17 6.72 0.33 ;
      RECT 6.13 0.17 6.22 0.33 ;
      RECT 4.5 0.19 4.95 0.28 ;
      RECT 7.63 0.17 7.72 0.355 ;
      RECT 5.22 0.17 7.72 0.26 ;
      RECT 5.33 0.625 5.42 0.965 ;
      RECT 4.61 0.625 4.7 0.95 ;
      RECT 4.61 0.625 7.855 0.715 ;
      RECT 5.4 0.35 5.49 0.715 ;
      RECT 4.68 0.37 4.77 0.715 ;
      RECT 1.82 0.665 1.91 1.15 ;
      RECT 1.32 0.665 1.41 1.15 ;
      RECT 0.82 0.665 0.91 1.15 ;
      RECT 0.32 0.665 0.41 1.15 ;
      RECT 0.07 0.665 2.16 0.755 ;
      RECT 2.07 0.37 2.16 0.755 ;
      RECT 2.07 0.625 4.145 0.715 ;
      RECT 1.57 0.37 1.66 0.755 ;
      RECT 1.07 0.37 1.16 0.755 ;
      RECT 0.57 0.27 0.66 0.755 ;
      RECT 0.07 0.255 0.16 0.755 ;
      RECT 7.785 1.08 9.855 1.17 ;
  END
END TINVX16H7R

MACRO TINVX1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TINVX1H7R 0 0 ;
  SIZE 1.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.2 1.48 ;
        RECT 0.31 1.075 0.45 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.2 0.08 ;
        RECT 0.295 -0.08 0.435 0.325 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.655 0.61 0.805 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.72 0.465 0.81 0.61 ;
        RECT 0.25 0.465 0.81 0.555 ;
        RECT 0.25 0.425 0.345 0.585 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.94 0.255 1.03 1.175 ;
        RECT 0.78 0.255 1.03 0.345 ;
      LAYER MET2 ;
        RECT 0.85 0.18 0.95 0.56 ;
      LAYER VIA1 ;
        RECT 0.855 0.255 0.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.07 0.225 0.16 1.135 ;
      RECT 0.07 0.895 0.85 0.985 ;
      RECT 0.76 0.72 0.85 0.985 ;
  END
END TINVX1H7R

MACRO TINVX1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TINVX1P4H7R 0 0 ;
  SIZE 1.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.4 1.48 ;
        RECT 0.295 1.095 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.4 0.08 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.641 0.575 0.821 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.695 0.455 0.785 0.625 ;
        RECT 0.225 0.455 0.785 0.545 ;
        RECT 0.225 0.455 0.315 0.625 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.795 1.095 1.185 1.185 ;
        RECT 1.095 0.255 1.185 1.185 ;
        RECT 0.795 0.255 1.185 0.345 ;
      LAYER MET2 ;
        RECT 1.05 0.18 1.15 0.56 ;
      LAYER VIA1 ;
        RECT 1.055 0.255 1.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.915 0.185 1.13 ;
      RECT 0.045 0.915 1.005 1.005 ;
      RECT 0.915 0.706 1.005 1.005 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 0.045 0.23 0.185 0.32 ;
  END
END TINVX1P4H7R

MACRO TINVX2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TINVX2H7R 0 0 ;
  SIZE 1.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 1.2 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 1.2 0.08 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.425 0.62 0.575 0.8 ;
      LAYER MET2 ;
        RECT 0.45 0.43 0.55 0.96 ;
      LAYER VIA1 ;
        RECT 0.455 0.655 0.545 0.745 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.525 0.17 1.1 0.26 ;
        RECT 0.225 0.415 0.615 0.505 ;
        RECT 0.525 0.17 0.615 0.505 ;
        RECT 0.225 0.415 0.345 0.575 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.04 0.825 1.145 1.17 ;
        RECT 1.055 0.375 1.145 1.17 ;
        RECT 0.76 0.375 1.145 0.465 ;
      LAYER MET2 ;
        RECT 1.05 0.625 1.15 1.16 ;
      LAYER VIA1 ;
        RECT 1.055 0.855 1.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.045 0.89 0.185 1.145 ;
      RECT 0.045 0.89 0.77 0.98 ;
      RECT 0.68 0.615 0.77 0.98 ;
      RECT 0.045 0.23 0.135 1.145 ;
      RECT 0.68 0.615 0.955 0.755 ;
      RECT 0.045 0.23 0.185 0.32 ;
  END
END TINVX2H7R

MACRO TINVX3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TINVX3H7R 0 0 ;
  SIZE 4.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.4 1.48 ;
        RECT 3.99 1.05 4.08 1.48 ;
        RECT 2.1 1.095 2.24 1.48 ;
        RECT 1.07 1.07 1.16 1.48 ;
        RECT 0.57 1.07 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.4 0.08 ;
        RECT 3.99 -0.08 4.08 0.33 ;
        RECT 3.49 -0.08 3.58 0.345 ;
        RECT 2.951 -0.08 3.091 0.305 ;
        RECT 1.335 -0.08 1.425 0.33 ;
        RECT 0.835 -0.08 0.925 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.25 0.425 0.565 0.575 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.395 0.625 1.575 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.24 0.205 4.33 1.04 ;
        RECT 3.74 0.855 4.33 0.945 ;
        RECT 3.904 0.42 4.33 0.51 ;
        RECT 3.83 0.401 3.942 0.459 ;
        RECT 3.786 0.368 3.904 0.414 ;
        RECT 3.876 0.42 4.33 0.496 ;
        RECT 3.74 0.331 3.876 0.369 ;
        RECT 3.74 0.855 3.83 1.04 ;
        RECT 3.74 0.205 3.83 0.369 ;
      LAYER MET2 ;
        RECT 4.05 0.63 4.15 1.16 ;
      LAYER VIA1 ;
        RECT 4.055 0.855 4.145 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.991 0.465 3.081 1.045 ;
      RECT 2.943 0.465 3.728 0.555 ;
      RECT 2.908 0.409 2.943 0.538 ;
      RECT 1.085 0.42 1.605 0.51 ;
      RECT 1.515 0.17 1.605 0.51 ;
      RECT 2.862 0.369 2.908 0.497 ;
      RECT 3.226 0.28 3.316 0.555 ;
      RECT 2.862 0.446 2.981 0.497 ;
      RECT 2.816 0.323 2.862 0.451 ;
      RECT 1.085 0.295 1.175 0.51 ;
      RECT 2.772 0.17 2.816 0.406 ;
      RECT 2.726 0.17 2.816 0.361 ;
      RECT 1.925 0.17 2.015 0.345 ;
      RECT 1.515 0.17 2.816 0.26 ;
      RECT 2.741 1.135 3.441 1.225 ;
      RECT 3.351 0.735 3.441 1.225 ;
      RECT 1.28 1.1 1.965 1.19 ;
      RECT 1.875 0.915 1.965 1.19 ;
      RECT 2.741 0.619 2.831 1.225 ;
      RECT 1.28 0.89 1.37 1.19 ;
      RECT 0.82 0.89 0.91 1.045 ;
      RECT 1.875 0.915 2.831 1.005 ;
      RECT 0.82 0.89 1.37 0.98 ;
      RECT 2.724 0.542 2.741 0.671 ;
      RECT 2.678 0.511 2.724 0.639 ;
      RECT 2.678 0.574 2.787 0.639 ;
      RECT 2.632 0.465 2.678 0.593 ;
      RECT 2.586 0.419 2.632 0.547 ;
      RECT 2.54 0.373 2.586 0.501 ;
      RECT 2.502 0.419 2.632 0.459 ;
      RECT 2.165 0.35 2.54 0.44 ;
      RECT 1.495 0.92 1.785 1.01 ;
      RECT 1.695 0.35 1.785 1.01 ;
      RECT 1.695 0.725 2.651 0.815 ;
      RECT 0.32 0.665 0.41 1.045 ;
      RECT 0.07 0.665 1.275 0.755 ;
      RECT 0.655 0.655 1.275 0.755 ;
      RECT 0.07 0.205 0.16 0.755 ;
      RECT 0.655 0.245 0.745 0.755 ;
      RECT 0.545 0.245 0.745 0.335 ;
  END
END TINVX3H7R

MACRO TINVX4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TINVX4H7R 0 0 ;
  SIZE 4.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.4 1.48 ;
        RECT 3.99 1.05 4.08 1.48 ;
        RECT 2.1 1.095 2.24 1.48 ;
        RECT 1.07 1.07 1.16 1.48 ;
        RECT 0.57 0.87 0.66 1.48 ;
        RECT 0.07 0.855 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.4 0.08 ;
        RECT 3.99 -0.08 4.08 0.33 ;
        RECT 3.49 -0.08 3.58 0.345 ;
        RECT 2.976 -0.08 3.066 0.33 ;
        RECT 1.335 -0.08 1.425 0.33 ;
        RECT 0.835 -0.08 0.925 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.455 0.565 0.555 ;
      LAYER MET2 ;
        RECT 0.25 0.225 0.35 0.76 ;
      LAYER VIA1 ;
        RECT 0.255 0.455 0.345 0.545 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.425 0.625 1.605 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.24 0.255 4.33 1.15 ;
        RECT 3.74 0.805 4.33 0.895 ;
        RECT 3.945 0.455 4.33 0.545 ;
        RECT 3.876 0.436 3.983 0.499 ;
        RECT 3.83 0.405 3.945 0.453 ;
        RECT 3.922 0.455 4.33 0.534 ;
        RECT 3.786 0.371 3.922 0.408 ;
        RECT 3.786 0.325 3.876 0.408 ;
        RECT 3.74 0.805 3.83 1.15 ;
        RECT 3.74 0.2 3.83 0.363 ;
      LAYER MET2 ;
        RECT 4.05 0.23 4.15 0.76 ;
      LAYER VIA1 ;
        RECT 4.055 0.455 4.145 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.991 0.465 3.081 0.95 ;
      RECT 2.943 0.465 3.73 0.555 ;
      RECT 2.908 0.409 2.943 0.538 ;
      RECT 1.085 0.42 1.605 0.51 ;
      RECT 1.515 0.17 1.605 0.51 ;
      RECT 2.862 0.369 2.908 0.497 ;
      RECT 3.226 0.355 3.316 0.555 ;
      RECT 2.862 0.446 2.981 0.497 ;
      RECT 2.816 0.323 2.862 0.451 ;
      RECT 1.085 0.37 1.175 0.51 ;
      RECT 2.772 0.17 2.816 0.406 ;
      RECT 2.726 0.17 2.816 0.361 ;
      RECT 1.925 0.17 2.015 0.355 ;
      RECT 1.515 0.17 2.816 0.26 ;
      RECT 0.82 0.87 0.91 1.21 ;
      RECT 1.28 1.1 1.965 1.19 ;
      RECT 1.875 0.85 1.965 1.19 ;
      RECT 2.541 1.075 3.556 1.165 ;
      RECT 3.216 0.875 3.556 1.165 ;
      RECT 1.28 0.87 1.37 1.19 ;
      RECT 2.541 0.85 2.831 1.165 ;
      RECT 2.741 0.549 2.831 1.165 ;
      RECT 0.82 0.87 1.37 0.96 ;
      RECT 1.875 0.85 2.831 0.94 ;
      RECT 2.701 0.461 2.741 0.589 ;
      RECT 2.701 0.504 2.787 0.589 ;
      RECT 2.655 0.418 2.701 0.546 ;
      RECT 2.617 0.395 2.655 0.504 ;
      RECT 2.15 0.395 2.655 0.485 ;
      RECT 1.495 0.92 1.785 1.01 ;
      RECT 1.695 0.35 1.785 1.01 ;
      RECT 1.695 0.635 2.62 0.725 ;
      RECT 0.32 0.665 0.41 1.15 ;
      RECT 0.045 0.665 1.275 0.755 ;
      RECT 0.655 0.255 0.745 0.755 ;
      RECT 0.045 0.24 0.135 0.755 ;
      RECT 0.545 0.255 0.745 0.345 ;
      RECT 0.045 0.24 0.185 0.33 ;
  END
END TINVX4H7R

MACRO TINVX6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TINVX6H7R 0 0 ;
  SIZE 5.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.6 1.48 ;
        RECT 5.19 1.07 5.28 1.48 ;
        RECT 4.69 1.055 4.78 1.48 ;
        RECT 2.71 1.07 2.8 1.48 ;
        RECT 2.105 1.225 2.245 1.48 ;
        RECT 1.32 1.055 1.41 1.48 ;
        RECT 0.795 0.895 0.935 1.48 ;
        RECT 0.295 0.895 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.6 0.08 ;
        RECT 5.305 -0.08 5.395 0.345 ;
        RECT 4.78 -0.08 4.92 0.305 ;
        RECT 4.285 -0.08 4.375 0.33 ;
        RECT 3.695 -0.08 3.835 0.175 ;
        RECT 2.065 -0.08 2.155 0.345 ;
        RECT 1.585 -0.08 1.675 0.33 ;
        RECT 1.085 -0.08 1.175 0.33 ;
        RECT 0.57 -0.08 0.66 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.405 0.515 0.745 0.605 ;
        RECT 0.655 0.425 0.745 0.605 ;
      LAYER MET2 ;
        RECT 0.65 0.225 0.75 0.76 ;
      LAYER VIA1 ;
        RECT 0.655 0.455 0.745 0.545 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.905 0.655 2.175 0.755 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.44 0.825 5.53 1.165 ;
        RECT 4.94 0.825 5.53 0.915 ;
        RECT 5.055 0.295 5.145 0.915 ;
        RECT 4.555 0.395 5.145 0.485 ;
        RECT 4.94 0.825 5.03 1.165 ;
        RECT 4.555 0.295 4.645 0.485 ;
      LAYER MET2 ;
        RECT 5.05 0.43 5.15 0.96 ;
      LAYER VIA1 ;
        RECT 5.055 0.655 5.145 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 3.63 1.08 4.435 1.17 ;
      RECT 3.63 1.08 4.481 1.147 ;
      RECT 4.397 1.061 4.527 1.101 ;
      RECT 4.435 1.019 4.527 1.101 ;
      RECT 4.435 1.019 4.573 1.055 ;
      RECT 4.481 0.973 4.595 1.021 ;
      RECT 4.527 0.927 4.641 0.987 ;
      RECT 4.573 0.893 4.595 1.021 ;
      RECT 4.595 0.575 4.685 0.942 ;
      RECT 4.035 0.575 4.685 0.665 ;
      RECT 4.035 0.265 4.125 0.665 ;
      RECT 1.335 0.435 2.335 0.525 ;
      RECT 2.245 0.175 2.335 0.525 ;
      RECT 1.835 0.355 1.925 0.525 ;
      RECT 1.335 0.36 1.425 0.525 ;
      RECT 3.405 0.265 4.125 0.355 ;
      RECT 2.905 0.175 2.995 0.33 ;
      RECT 2.245 0.175 3.495 0.265 ;
      RECT 2.96 1.12 3.495 1.21 ;
      RECT 3.405 0.87 3.495 1.21 ;
      RECT 1.57 0.855 1.66 1.195 ;
      RECT 1.07 0.855 1.16 1.195 ;
      RECT 1.57 1.03 2.55 1.12 ;
      RECT 2.46 0.87 2.55 1.12 ;
      RECT 2.96 0.87 3.05 1.21 ;
      RECT 3.405 0.87 3.995 0.96 ;
      RECT 3.855 0.773 3.995 0.96 ;
      RECT 2.46 0.87 3.05 0.96 ;
      RECT 1.07 0.855 1.66 0.945 ;
      RECT 3.855 0.773 4.48 0.863 ;
      RECT 3.855 0.445 3.945 0.96 ;
      RECT 2.655 0.445 3.945 0.535 ;
      RECT 3.155 0.37 3.245 0.535 ;
      RECT 2.655 0.355 2.745 0.535 ;
      RECT 1.775 0.85 2.37 0.94 ;
      RECT 2.28 0.665 2.37 0.94 ;
      RECT 2.28 0.665 3.7 0.755 ;
      RECT 2.425 0.355 2.515 0.755 ;
      RECT 0.07 0.545 0.16 1.165 ;
      RECT 0.57 0.7 0.66 1.15 ;
      RECT 0.07 0.7 0.91 0.79 ;
      RECT 0.835 0.665 1.67 0.755 ;
      RECT 0.835 0.22 0.925 0.755 ;
      RECT 0.116 0.5 0.206 0.583 ;
      RECT 0.16 0.455 0.252 0.537 ;
      RECT 0.16 0.455 0.298 0.491 ;
      RECT 0.206 0.409 0.32 0.457 ;
      RECT 0.252 0.363 0.366 0.423 ;
      RECT 0.298 0.329 0.32 0.457 ;
      RECT 0.32 0.215 0.41 0.378 ;
  END
END TINVX6H7R

MACRO TINVX8H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TINVX8H7R 0 0 ;
  SIZE 7.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 7.2 1.48 ;
        RECT 6.691 1.095 6.831 1.48 ;
        RECT 6.191 1.095 6.331 1.48 ;
        RECT 5.716 1.055 5.806 1.48 ;
        RECT 4.102 1.205 4.242 1.48 ;
        RECT 3.562 1.07 3.652 1.48 ;
        RECT 2.997 1.2 3.087 1.48 ;
        RECT 2.07 1.07 2.16 1.48 ;
        RECT 1.57 1.07 1.66 1.48 ;
        RECT 1.07 0.87 1.16 1.48 ;
        RECT 0.57 0.87 0.66 1.48 ;
        RECT 0.07 0.855 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 7.2 0.08 ;
        RECT 7.022 -0.08 7.112 0.345 ;
        RECT 6.491 -0.08 6.631 0.305 ;
        RECT 5.991 -0.08 6.131 0.305 ;
        RECT 5.261 -0.08 5.401 0.305 ;
        RECT 4.761 -0.08 4.901 0.305 ;
        RECT 3.29 -0.08 3.38 0.33 ;
        RECT 2.57 -0.08 2.66 0.33 ;
        RECT 2.045 -0.08 2.185 0.305 ;
        RECT 1.57 -0.08 1.66 0.33 ;
        RECT 1.07 -0.08 1.16 0.33 ;
        RECT 0.57 -0.08 0.66 0.33 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1 0.435 1.225 0.555 ;
      LAYER MET2 ;
        RECT 1.05 0.225 1.15 0.76 ;
      LAYER VIA1 ;
        RECT 1.055 0.455 1.145 0.545 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.57 0.65 2.84 0.75 ;
      LAYER MET2 ;
        RECT 2.65 0.43 2.75 0.96 ;
      LAYER VIA1 ;
        RECT 2.655 0.655 2.745 0.745 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.966 0.855 7.056 1.041 ;
        RECT 6.766 0.855 7.056 1.005 ;
        RECT 6.766 0.31 6.856 1.005 ;
        RECT 6.012 0.934 7.056 1.005 ;
        RECT 6.05 0.915 7.056 1.005 ;
        RECT 5.766 0.395 6.856 0.485 ;
        RECT 6.266 0.31 6.356 0.485 ;
        RECT 5.966 0.976 6.088 1.021 ;
        RECT 5.966 0.976 6.056 1.139 ;
        RECT 5.766 0.295 5.856 0.485 ;
      LAYER MET2 ;
        RECT 6.85 0.63 6.95 1.16 ;
      LAYER VIA1 ;
        RECT 6.855 0.855 6.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 3.812 0.87 3.902 1.21 ;
      RECT 3.312 0.87 3.402 1.21 ;
      RECT 1.82 0.87 1.91 1.21 ;
      RECT 1.32 0.87 1.41 1.21 ;
      RECT 2.347 1.114 2.862 1.204 ;
      RECT 2.347 1.114 2.908 1.181 ;
      RECT 3.812 1.025 5.576 1.115 ;
      RECT 5.486 0.867 5.576 1.115 ;
      RECT 2.824 1.095 2.956 1.129 ;
      RECT 2.908 1.025 2.918 1.153 ;
      RECT 2.347 0.87 2.437 1.204 ;
      RECT 2.918 1.02 3.402 1.11 ;
      RECT 2.862 1.053 3.402 1.11 ;
      RECT 4.505 0.6 4.595 1.115 ;
      RECT 3.312 0.87 3.902 0.96 ;
      RECT 1.32 0.87 2.437 0.96 ;
      RECT 5.486 0.867 5.727 0.957 ;
      RECT 5.486 0.867 5.773 0.934 ;
      RECT 5.689 0.848 5.815 0.89 ;
      RECT 5.727 0.806 5.853 0.85 ;
      RECT 5.773 0.762 5.815 0.89 ;
      RECT 5.815 0.741 6.011 0.831 ;
      RECT 4.286 0.6 4.595 0.69 ;
      RECT 4.286 0.37 4.376 0.69 ;
      RECT 3.761 0.42 4.376 0.51 ;
      RECT 3.761 0.355 3.901 0.51 ;
      RECT 4.711 0.845 5.351 0.935 ;
      RECT 5.036 0.395 5.126 0.935 ;
      RECT 5.536 0.59 5.731 0.68 ;
      RECT 5.536 0.242 5.626 0.68 ;
      RECT 3.11 0.42 3.626 0.51 ;
      RECT 3.536 0.17 3.626 0.51 ;
      RECT 2.415 0.42 2.84 0.51 ;
      RECT 2.75 0.17 2.84 0.51 ;
      RECT 4.536 0.395 5.626 0.485 ;
      RECT 1.795 0.395 2.505 0.485 ;
      RECT 3.11 0.17 3.2 0.51 ;
      RECT 4.536 0.17 4.626 0.485 ;
      RECT 4.036 0.17 4.126 0.33 ;
      RECT 3.536 0.17 4.626 0.26 ;
      RECT 2.75 0.17 3.2 0.26 ;
      RECT 2.682 0.84 2.772 1.02 ;
      RECT 2.682 0.84 3.02 0.93 ;
      RECT 2.93 0.37 3.02 0.93 ;
      RECT 4.082 0.812 4.415 0.902 ;
      RECT 4.082 0.69 4.172 0.902 ;
      RECT 2.93 0.69 4.172 0.78 ;
      RECT 0.82 0.27 0.91 1.15 ;
      RECT 0.32 0.27 0.41 1.15 ;
      RECT 0.32 0.645 1.95 0.735 ;
      RECT 1.32 0.27 1.41 0.735 ;
  END
END TINVX8H7R

MACRO XNOR2X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2X0P5H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.575 1.2 1.665 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.59 -0.08 1.68 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.505 1.555 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.795 0.405 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.84 0.205 1.945 1.175 ;
      LAYER MET2 ;
        RECT 1.85 0.84 1.95 1.22 ;
      LAYER VIA1 ;
        RECT 1.855 1.055 1.945 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.78 1.11 1.446 1.2 ;
      RECT 0.78 1.11 1.492 1.177 ;
      RECT 1.408 1.091 1.538 1.131 ;
      RECT 0.78 0.35 0.87 1.2 ;
      RECT 1.446 1.049 1.538 1.131 ;
      RECT 1.492 1.003 1.584 1.085 ;
      RECT 1.492 1.003 1.63 1.039 ;
      RECT 1.538 0.957 1.65 1.006 ;
      RECT 1.584 0.911 1.696 0.973 ;
      RECT 1.63 0.878 1.65 1.006 ;
      RECT 1.65 0.766 1.74 0.928 ;
      RECT 0.78 0.35 0.925 0.44 ;
      RECT 1.275 0.744 1.365 1.018 ;
      RECT 1.246 0.744 1.365 0.783 ;
      RECT 1.2 0.468 1.29 0.745 ;
      RECT 1.2 0.707 1.336 0.745 ;
      RECT 1.2 0.468 1.336 0.506 ;
      RECT 1.246 0.43 1.34 0.481 ;
      RECT 1.275 0.408 1.386 0.456 ;
      RECT 1.336 0.353 1.34 0.481 ;
      RECT 1.34 0.205 1.43 0.411 ;
      RECT 1.29 0.378 1.43 0.411 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 1.02 0.84 1.16 0.93 ;
      RECT 1.02 0.17 1.11 0.93 ;
      RECT 0.045 0.445 0.64 0.535 ;
      RECT 0.55 0.17 0.64 0.535 ;
      RECT 1.02 0.17 1.18 0.345 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.55 0.17 1.18 0.26 ;
  END
END XNOR2X0P5H7R

MACRO XNOR2X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2X0P7H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.575 1.2 1.665 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.59 -0.08 1.68 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.475 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.795 0.405 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.84 0.225 1.945 1.103 ;
      LAYER MET2 ;
        RECT 1.85 0.18 1.95 0.56 ;
      LAYER VIA1 ;
        RECT 1.855 0.255 1.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.78 1.11 1.446 1.2 ;
      RECT 0.78 1.11 1.492 1.177 ;
      RECT 1.408 1.091 1.538 1.131 ;
      RECT 0.78 0.35 0.87 1.2 ;
      RECT 1.446 1.049 1.538 1.131 ;
      RECT 1.492 1.003 1.584 1.085 ;
      RECT 1.492 1.003 1.63 1.039 ;
      RECT 1.538 0.957 1.65 1.006 ;
      RECT 1.584 0.911 1.696 0.973 ;
      RECT 1.63 0.878 1.65 1.006 ;
      RECT 1.65 0.753 1.74 0.928 ;
      RECT 0.78 0.35 0.925 0.44 ;
      RECT 1.275 0.732 1.365 1.018 ;
      RECT 1.241 0.692 1.331 0.77 ;
      RECT 1.195 0.453 1.285 0.73 ;
      RECT 1.195 0.453 1.331 0.491 ;
      RECT 1.241 0.413 1.34 0.464 ;
      RECT 1.275 0.391 1.386 0.436 ;
      RECT 1.331 0.335 1.34 0.464 ;
      RECT 1.34 0.205 1.43 0.391 ;
      RECT 1.285 0.363 1.43 0.391 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 1.015 0.84 1.16 0.93 ;
      RECT 1.015 0.17 1.105 0.93 ;
      RECT 0.045 0.445 0.64 0.535 ;
      RECT 0.55 0.17 0.64 0.535 ;
      RECT 1.015 0.17 1.18 0.345 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.55 0.17 1.18 0.26 ;
  END
END XNOR2X0P7H7R

MACRO XNOR2X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2X1H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.575 1.2 1.665 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.565 -0.08 1.705 0.305 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.475 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.795 0.405 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.84 0.225 1.945 1.055 ;
      LAYER MET2 ;
        RECT 1.85 0.18 1.95 0.56 ;
      LAYER VIA1 ;
        RECT 1.855 0.255 1.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.78 1.11 1.446 1.2 ;
      RECT 0.78 1.11 1.492 1.177 ;
      RECT 1.408 1.091 1.538 1.131 ;
      RECT 0.78 0.35 0.87 1.2 ;
      RECT 1.446 1.049 1.538 1.131 ;
      RECT 1.492 1.003 1.584 1.085 ;
      RECT 1.492 1.003 1.63 1.039 ;
      RECT 1.538 0.957 1.65 1.006 ;
      RECT 1.584 0.911 1.696 0.973 ;
      RECT 1.63 0.878 1.65 1.006 ;
      RECT 1.65 0.73 1.74 0.928 ;
      RECT 0.78 0.35 0.925 0.44 ;
      RECT 1.275 0.747 1.365 1.018 ;
      RECT 1.241 0.707 1.331 0.785 ;
      RECT 1.195 0.453 1.285 0.745 ;
      RECT 1.195 0.453 1.331 0.491 ;
      RECT 1.241 0.413 1.34 0.464 ;
      RECT 1.275 0.391 1.386 0.436 ;
      RECT 1.331 0.335 1.34 0.464 ;
      RECT 1.34 0.205 1.43 0.391 ;
      RECT 1.285 0.363 1.43 0.391 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 1.015 0.865 1.16 0.955 ;
      RECT 1.015 0.17 1.105 0.955 ;
      RECT 0.045 0.445 0.64 0.535 ;
      RECT 0.55 0.17 0.64 0.535 ;
      RECT 1.015 0.17 1.18 0.345 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.55 0.17 1.18 0.26 ;
  END
END XNOR2X1H7R

MACRO XNOR2X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2X1P4H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.575 1.2 1.665 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.59 -0.08 1.68 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.475 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.345 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.84 0.916 1.955 1.056 ;
        RECT 1.865 0.301 1.955 1.056 ;
        RECT 1.84 0.301 1.955 0.575 ;
      LAYER MET2 ;
        RECT 1.85 0.225 1.95 0.76 ;
      LAYER VIA1 ;
        RECT 1.855 0.455 1.945 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.78 1.14 1.394 1.23 ;
      RECT 0.78 1.14 1.44 1.207 ;
      RECT 1.356 1.121 1.486 1.161 ;
      RECT 0.78 0.35 0.87 1.23 ;
      RECT 1.394 1.079 1.486 1.161 ;
      RECT 1.44 1.033 1.532 1.115 ;
      RECT 1.486 0.987 1.578 1.069 ;
      RECT 1.532 0.941 1.624 1.023 ;
      RECT 1.532 0.941 1.67 0.977 ;
      RECT 1.578 0.895 1.685 0.947 ;
      RECT 1.624 0.849 1.731 0.916 ;
      RECT 1.67 0.818 1.685 0.947 ;
      RECT 1.685 0.66 1.775 0.871 ;
      RECT 0.78 0.35 0.925 0.44 ;
      RECT 1.275 0.712 1.365 0.998 ;
      RECT 1.241 0.672 1.331 0.75 ;
      RECT 1.195 0.438 1.285 0.71 ;
      RECT 1.195 0.438 1.331 0.476 ;
      RECT 1.241 0.398 1.34 0.449 ;
      RECT 1.275 0.376 1.386 0.421 ;
      RECT 1.331 0.32 1.34 0.449 ;
      RECT 1.34 0.205 1.43 0.376 ;
      RECT 1.285 0.348 1.43 0.376 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 1.015 0.865 1.16 0.955 ;
      RECT 1.015 0.17 1.105 0.955 ;
      RECT 0.045 0.445 0.64 0.535 ;
      RECT 0.55 0.17 0.64 0.535 ;
      RECT 1.015 0.17 1.18 0.345 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.55 0.17 1.18 0.26 ;
  END
END XNOR2X1P4H7R

MACRO XNOR2X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2X2H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 2.09 1.035 2.18 1.48 ;
        RECT 1.575 1.2 1.665 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 2.09 -0.08 2.18 0.345 ;
        RECT 1.59 -0.08 1.68 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.5 1.545 0.8 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.345 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.815 1.005 2 1.095 ;
        RECT 1.91 0.245 2 1.095 ;
        RECT 1.815 0.245 2 0.345 ;
      LAYER MET2 ;
        RECT 1.85 0.18 1.95 0.56 ;
      LAYER VIA1 ;
        RECT 1.855 0.255 1.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.78 1.14 1.416 1.23 ;
      RECT 0.78 1.14 1.462 1.207 ;
      RECT 1.378 1.121 1.508 1.161 ;
      RECT 0.78 0.35 0.87 1.23 ;
      RECT 1.416 1.079 1.508 1.161 ;
      RECT 1.462 1.033 1.554 1.115 ;
      RECT 1.508 0.987 1.6 1.069 ;
      RECT 1.554 0.941 1.646 1.023 ;
      RECT 1.6 0.895 1.692 0.977 ;
      RECT 1.646 0.849 1.766 0.898 ;
      RECT 1.692 0.807 1.73 0.935 ;
      RECT 1.73 0.686 1.82 0.88 ;
      RECT 0.78 0.35 0.93 0.44 ;
      RECT 1.275 0.793 1.365 1.018 ;
      RECT 1.246 0.793 1.365 0.832 ;
      RECT 1.2 0.443 1.29 0.794 ;
      RECT 1.2 0.756 1.336 0.794 ;
      RECT 1.2 0.443 1.336 0.481 ;
      RECT 1.246 0.405 1.34 0.456 ;
      RECT 1.275 0.383 1.386 0.431 ;
      RECT 1.336 0.328 1.34 0.456 ;
      RECT 1.34 0.205 1.43 0.386 ;
      RECT 1.29 0.353 1.43 0.386 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 1.02 0.865 1.16 0.955 ;
      RECT 1.02 0.17 1.11 0.955 ;
      RECT 0.045 0.445 0.64 0.535 ;
      RECT 0.55 0.17 0.64 0.535 ;
      RECT 1.02 0.17 1.185 0.345 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.55 0.17 1.185 0.26 ;
  END
END XNOR2X2H7R

MACRO XNOR2X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2X3H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 2.09 1.035 2.18 1.48 ;
        RECT 1.575 1.2 1.665 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 2.09 -0.08 2.18 0.345 ;
        RECT 1.59 -0.08 1.68 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.475 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.235 0.74 0.35 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.815 0.97 2 1.06 ;
        RECT 1.91 0.255 2 1.06 ;
        RECT 1.815 0.255 2 0.345 ;
      LAYER MET2 ;
        RECT 1.85 0.18 1.95 0.56 ;
      LAYER VIA1 ;
        RECT 1.855 0.255 1.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.78 1.14 1.416 1.23 ;
      RECT 0.78 1.14 1.462 1.207 ;
      RECT 1.378 1.121 1.508 1.161 ;
      RECT 0.78 0.35 0.87 1.23 ;
      RECT 1.416 1.079 1.508 1.161 ;
      RECT 1.462 1.033 1.554 1.115 ;
      RECT 1.508 0.987 1.6 1.069 ;
      RECT 1.554 0.941 1.646 1.023 ;
      RECT 1.6 0.895 1.692 0.977 ;
      RECT 1.646 0.849 1.766 0.898 ;
      RECT 1.692 0.807 1.73 0.935 ;
      RECT 1.73 0.715 1.82 0.88 ;
      RECT 0.78 0.35 0.93 0.44 ;
      RECT 1.275 0.793 1.365 1.018 ;
      RECT 1.246 0.793 1.365 0.832 ;
      RECT 1.2 0.438 1.29 0.794 ;
      RECT 1.2 0.756 1.336 0.794 ;
      RECT 1.2 0.438 1.336 0.476 ;
      RECT 1.246 0.4 1.34 0.451 ;
      RECT 1.275 0.378 1.386 0.426 ;
      RECT 1.336 0.323 1.34 0.451 ;
      RECT 1.34 0.205 1.43 0.381 ;
      RECT 1.29 0.348 1.43 0.381 ;
      RECT 0.045 1.05 0.185 1.14 ;
      RECT 0.045 0.23 0.135 1.14 ;
      RECT 1.02 0.865 1.16 0.955 ;
      RECT 1.02 0.17 1.11 0.955 ;
      RECT 0.045 0.49 0.64 0.58 ;
      RECT 0.55 0.17 0.64 0.58 ;
      RECT 1.02 0.17 1.185 0.345 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.55 0.17 1.185 0.26 ;
  END
END XNOR2X3H7R

MACRO XNOR2X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2X4H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 2.09 1.035 2.18 1.48 ;
        RECT 1.575 1.2 1.665 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 2.083 -0.08 2.223 0.305 ;
        RECT 1.605 -0.08 1.695 0.33 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.52 1.545 0.82 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.855 0.395 2.448 0.485 ;
        RECT 2.358 0.255 2.448 0.485 ;
        RECT 1.815 0.97 2 1.06 ;
        RECT 1.91 0.395 2 1.06 ;
        RECT 1.855 0.225 1.945 0.485 ;
      LAYER MET2 ;
        RECT 1.85 0.18 1.95 0.56 ;
      LAYER VIA1 ;
        RECT 1.855 0.255 1.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.78 1.14 1.416 1.23 ;
      RECT 0.78 1.14 1.462 1.207 ;
      RECT 1.378 1.121 1.508 1.161 ;
      RECT 0.78 0.35 0.87 1.23 ;
      RECT 1.416 1.079 1.508 1.161 ;
      RECT 1.462 1.033 1.554 1.115 ;
      RECT 1.508 0.987 1.6 1.069 ;
      RECT 1.554 0.941 1.646 1.023 ;
      RECT 1.6 0.895 1.692 0.977 ;
      RECT 1.646 0.849 1.766 0.898 ;
      RECT 1.692 0.807 1.73 0.935 ;
      RECT 1.73 0.62 1.82 0.88 ;
      RECT 0.78 0.35 0.93 0.44 ;
      RECT 1.275 0.797 1.365 1.005 ;
      RECT 1.254 0.797 1.365 0.836 ;
      RECT 1.208 0.475 1.298 0.802 ;
      RECT 1.208 0.764 1.344 0.802 ;
      RECT 1.208 0.475 1.344 0.513 ;
      RECT 1.254 0.441 1.355 0.485 ;
      RECT 1.275 0.419 1.401 0.456 ;
      RECT 1.344 0.356 1.355 0.485 ;
      RECT 1.298 0.385 1.401 0.456 ;
      RECT 1.355 0.225 1.445 0.411 ;
      RECT 0.07 0.89 0.16 1.035 ;
      RECT 0.07 0.89 0.51 0.98 ;
      RECT 0.42 0.395 0.51 0.98 ;
      RECT 1.02 0.865 1.16 0.955 ;
      RECT 1.02 0.17 1.11 0.955 ;
      RECT 0.07 0.395 0.64 0.485 ;
      RECT 0.55 0.17 0.64 0.485 ;
      RECT 0.07 0.305 0.16 0.485 ;
      RECT 1.02 0.17 1.215 0.345 ;
      RECT 0.55 0.17 1.215 0.26 ;
  END
END XNOR2X4H7R

MACRO XNOR2X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2X6H7R 0 0 ;
  SIZE 3.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3.2 1.48 ;
        RECT 2.368 1.05 2.458 1.48 ;
        RECT 1.853 1.2 1.943 1.48 ;
        RECT 0.57 1.07 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3.2 0.08 ;
        RECT 2.868 -0.08 2.958 0.345 ;
        RECT 2.343 -0.08 2.483 0.305 ;
        RECT 1.868 -0.08 1.958 0.33 ;
        RECT 0.545 -0.08 0.685 0.305 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.73 0.51 1.945 0.6 ;
        RECT 1.855 0.425 1.945 0.6 ;
      LAYER MET2 ;
        RECT 1.85 0.225 1.95 0.76 ;
      LAYER VIA1 ;
        RECT 1.855 0.455 1.945 0.545 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.195 0.655 0.535 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.618 0.295 2.708 0.945 ;
        RECT 2.164 0.872 2.708 0.945 ;
        RECT 2.199 0.855 2.708 0.945 ;
        RECT 2.118 0.395 2.708 0.485 ;
        RECT 2.118 0.913 2.237 0.96 ;
        RECT 2.118 0.913 2.208 1.08 ;
        RECT 2.118 0.295 2.208 0.485 ;
      LAYER MET2 ;
        RECT 2.45 0.625 2.55 1.16 ;
      LAYER VIA1 ;
        RECT 2.455 0.855 2.545 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.03 1.11 1.701 1.2 ;
      RECT 1.03 1.11 1.747 1.177 ;
      RECT 1.663 1.091 1.793 1.131 ;
      RECT 1.03 0.35 1.12 1.2 ;
      RECT 1.701 1.049 1.793 1.131 ;
      RECT 1.747 1.003 1.839 1.085 ;
      RECT 1.793 0.957 1.885 1.039 ;
      RECT 1.839 0.911 1.931 0.993 ;
      RECT 1.885 0.865 1.977 0.947 ;
      RECT 1.931 0.819 2.023 0.901 ;
      RECT 1.977 0.773 2.069 0.855 ;
      RECT 1.977 0.773 2.115 0.809 ;
      RECT 2.023 0.727 2.128 0.78 ;
      RECT 2.023 0.727 2.166 0.754 ;
      RECT 2.128 0.645 2.468 0.735 ;
      RECT 2.069 0.681 2.468 0.735 ;
      RECT 2.115 0.651 2.128 0.78 ;
      RECT 1.03 0.35 1.175 0.44 ;
      RECT 1.525 0.762 1.615 1.018 ;
      RECT 1.514 0.762 1.615 0.801 ;
      RECT 1.468 0.485 1.558 0.772 ;
      RECT 1.468 0.734 1.604 0.772 ;
      RECT 1.468 0.485 1.604 0.523 ;
      RECT 1.514 0.456 1.618 0.493 ;
      RECT 1.525 0.434 1.664 0.463 ;
      RECT 1.604 0.365 1.618 0.493 ;
      RECT 1.558 0.395 1.664 0.463 ;
      RECT 1.618 0.255 1.708 0.418 ;
      RECT 0.32 0.89 0.41 1.14 ;
      RECT 0.32 0.89 0.76 0.98 ;
      RECT 0.67 0.395 0.76 0.98 ;
      RECT 1.27 0.82 1.41 0.91 ;
      RECT 1.27 0.17 1.36 0.91 ;
      RECT 0.32 0.395 0.89 0.485 ;
      RECT 0.8 0.17 0.89 0.485 ;
      RECT 0.32 0.22 0.41 0.485 ;
      RECT 1.27 0.17 1.478 0.35 ;
      RECT 0.8 0.17 1.478 0.26 ;
  END
END XNOR2X6H7R

MACRO XNOR3X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR3X0P5H7R 0 0 ;
  SIZE 4.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.2 1.48 ;
        RECT 3.29 1.05 3.38 1.48 ;
        RECT 2.81 1.035 2.9 1.48 ;
        RECT 1.575 1.2 1.665 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.2 0.08 ;
        RECT 3.76 -0.08 3.85 0.33 ;
        RECT 3.28 -0.08 3.37 0.345 ;
        RECT 1.59 -0.08 1.68 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.51 1.555 0.78 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.345 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.22 0.81 3.42 0.945 ;
      LAYER MET2 ;
        RECT 3.25 0.63 3.35 1.16 ;
      LAYER VIA1 ;
        RECT 3.255 0.855 3.345 0.945 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.68 1.055 4.1 1.145 ;
        RECT 4.01 0.205 4.1 1.145 ;
      LAYER MET2 ;
        RECT 3.85 0.84 3.95 1.22 ;
      LAYER VIA1 ;
        RECT 3.855 1.055 3.945 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.335 0.435 2.425 1.015 ;
      RECT 3.83 0.62 3.92 0.76 ;
      RECT 2.335 0.62 3.92 0.71 ;
      RECT 2.07 0.435 2.665 0.525 ;
      RECT 2.525 0.35 2.665 0.525 ;
      RECT 2.07 0.205 2.16 0.525 ;
      RECT 2.775 0.44 3.6 0.53 ;
      RECT 3.51 0.205 3.6 0.53 ;
      RECT 2.775 0.35 2.915 0.53 ;
      RECT 2.07 1.14 2.72 1.23 ;
      RECT 2.63 0.835 2.72 1.23 ;
      RECT 2.07 1.035 2.16 1.23 ;
      RECT 3.04 0.967 3.13 1.135 ;
      RECT 3.022 0.89 3.04 1.018 ;
      RECT 2.976 0.858 3.022 0.986 ;
      RECT 2.976 0.922 3.086 0.986 ;
      RECT 2.938 0.922 3.086 0.944 ;
      RECT 2.63 0.835 2.976 0.925 ;
      RECT 3.03 0.17 3.12 0.345 ;
      RECT 2.32 0.17 2.41 0.345 ;
      RECT 2.32 0.17 3.12 0.26 ;
      RECT 1.84 0.205 1.93 1.135 ;
      RECT 1.84 0.669 2.01 0.809 ;
      RECT 0.78 1.14 1.416 1.23 ;
      RECT 0.78 1.14 1.462 1.207 ;
      RECT 1.378 1.121 1.508 1.161 ;
      RECT 0.78 0.43 0.87 1.23 ;
      RECT 1.416 1.079 1.508 1.161 ;
      RECT 1.462 1.033 1.554 1.115 ;
      RECT 1.508 0.987 1.6 1.069 ;
      RECT 1.508 0.987 1.646 1.023 ;
      RECT 1.554 0.941 1.65 0.998 ;
      RECT 1.6 0.895 1.696 0.973 ;
      RECT 1.646 0.87 1.65 0.998 ;
      RECT 1.65 0.765 1.74 0.928 ;
      RECT 0.78 0.43 0.92 0.52 ;
      RECT 1.275 0.823 1.365 1.018 ;
      RECT 1.24 0.438 1.33 0.862 ;
      RECT 1.225 0.635 1.33 0.837 ;
      RECT 1.275 0.398 1.386 0.461 ;
      RECT 1.33 0.361 1.34 0.489 ;
      RECT 1.34 0.205 1.43 0.416 ;
      RECT 1.321 0.37 1.43 0.416 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 1.02 0.96 1.16 1.05 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 1.02 0.25 1.11 1.05 ;
      RECT 1.02 0.405 1.15 0.545 ;
      RECT 0.045 0.445 0.64 0.535 ;
      RECT 0.55 0.25 0.64 0.535 ;
      RECT 0.55 0.25 1.11 0.34 ;
      RECT 0.045 0.23 0.185 0.32 ;
  END
END XNOR3X0P5H7R

MACRO XNOR3X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR3X0P7H7R 0 0 ;
  SIZE 4.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.2 1.48 ;
        RECT 3.29 1.05 3.38 1.48 ;
        RECT 2.81 1.035 2.9 1.48 ;
        RECT 1.575 1.2 1.665 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.2 0.08 ;
        RECT 3.76 -0.08 3.85 0.33 ;
        RECT 3.28 -0.08 3.37 0.345 ;
        RECT 1.59 -0.08 1.68 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.51 1.555 0.78 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.345 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.22 0.8 3.4 0.95 ;
      LAYER MET2 ;
        RECT 3.25 0.63 3.35 1.16 ;
      LAYER VIA1 ;
        RECT 3.255 0.855 3.345 0.945 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.68 1.055 4.1 1.145 ;
        RECT 4.01 0.229 4.1 1.145 ;
      LAYER MET2 ;
        RECT 3.85 0.84 3.95 1.22 ;
      LAYER VIA1 ;
        RECT 3.855 1.055 3.945 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.335 0.435 2.425 1.015 ;
      RECT 3.83 0.62 3.92 0.76 ;
      RECT 2.335 0.62 3.92 0.71 ;
      RECT 2.07 0.435 2.665 0.525 ;
      RECT 2.525 0.35 2.665 0.525 ;
      RECT 2.07 0.205 2.16 0.525 ;
      RECT 2.775 0.44 3.6 0.53 ;
      RECT 3.51 0.205 3.6 0.53 ;
      RECT 2.775 0.35 2.915 0.53 ;
      RECT 2.07 1.105 2.72 1.195 ;
      RECT 2.63 0.835 2.72 1.195 ;
      RECT 3.04 0.967 3.13 1.135 ;
      RECT 2.07 1.035 2.16 1.195 ;
      RECT 3.022 0.89 3.04 1.018 ;
      RECT 2.976 0.858 3.022 0.986 ;
      RECT 2.976 0.922 3.086 0.986 ;
      RECT 2.938 0.922 3.086 0.944 ;
      RECT 2.63 0.835 2.976 0.925 ;
      RECT 3.03 0.17 3.12 0.345 ;
      RECT 2.32 0.17 2.41 0.345 ;
      RECT 2.32 0.17 3.12 0.26 ;
      RECT 1.84 0.205 1.93 1.135 ;
      RECT 1.84 0.669 2.01 0.809 ;
      RECT 0.78 1.14 1.416 1.23 ;
      RECT 0.78 1.14 1.462 1.207 ;
      RECT 1.378 1.121 1.508 1.161 ;
      RECT 0.78 0.43 0.87 1.23 ;
      RECT 1.416 1.079 1.508 1.161 ;
      RECT 1.462 1.033 1.554 1.115 ;
      RECT 1.508 0.987 1.6 1.069 ;
      RECT 1.508 0.987 1.646 1.023 ;
      RECT 1.554 0.941 1.65 0.998 ;
      RECT 1.6 0.895 1.696 0.973 ;
      RECT 1.646 0.87 1.65 0.998 ;
      RECT 1.65 0.765 1.74 0.928 ;
      RECT 0.78 0.43 0.92 0.52 ;
      RECT 1.275 0.823 1.365 1.018 ;
      RECT 1.24 0.408 1.33 0.862 ;
      RECT 1.225 0.635 1.33 0.837 ;
      RECT 1.275 0.368 1.386 0.431 ;
      RECT 1.33 0.331 1.34 0.459 ;
      RECT 1.34 0.205 1.43 0.386 ;
      RECT 1.321 0.34 1.43 0.386 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 1.02 0.96 1.16 1.05 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 1.02 0.17 1.11 1.05 ;
      RECT 1.02 0.405 1.15 0.545 ;
      RECT 0.045 0.445 0.64 0.535 ;
      RECT 0.55 0.17 0.64 0.535 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.55 0.17 1.11 0.26 ;
  END
END XNOR3X0P7H7R

MACRO XNOR3X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR3X1H7R 0 0 ;
  SIZE 4.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.2 1.48 ;
        RECT 3.29 1.05 3.38 1.48 ;
        RECT 2.81 1.035 2.9 1.48 ;
        RECT 1.575 1.2 1.665 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.2 0.08 ;
        RECT 3.76 -0.08 3.85 0.33 ;
        RECT 3.28 -0.08 3.37 0.345 ;
        RECT 1.59 -0.08 1.68 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.505 1.555 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.345 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.35 0.655 3.65 0.745 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.68 1.055 4.1 1.145 ;
        RECT 4.01 0.265 4.1 1.145 ;
      LAYER MET2 ;
        RECT 3.85 0.84 3.95 1.22 ;
      LAYER VIA1 ;
        RECT 3.855 1.055 3.945 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.335 0.435 2.425 1.015 ;
      RECT 3.214 0.855 3.92 0.945 ;
      RECT 3.83 0.705 3.92 0.945 ;
      RECT 3.201 0.81 3.214 0.939 ;
      RECT 3.155 0.781 3.201 0.909 ;
      RECT 3.109 0.735 3.155 0.863 ;
      RECT 3.109 0.836 3.252 0.863 ;
      RECT 3.063 0.689 3.109 0.817 ;
      RECT 3.017 0.643 3.063 0.771 ;
      RECT 2.979 0.689 3.109 0.729 ;
      RECT 2.335 0.62 3.017 0.71 ;
      RECT 2.07 0.435 2.665 0.525 ;
      RECT 2.525 0.35 2.665 0.525 ;
      RECT 2.07 0.205 2.16 0.525 ;
      RECT 2.775 0.44 3.6 0.53 ;
      RECT 3.51 0.205 3.6 0.53 ;
      RECT 2.775 0.35 2.915 0.53 ;
      RECT 2.07 1.105 2.72 1.195 ;
      RECT 2.63 0.835 2.72 1.195 ;
      RECT 3.04 0.967 3.13 1.135 ;
      RECT 2.07 1.035 2.16 1.195 ;
      RECT 3.022 0.89 3.04 1.018 ;
      RECT 2.976 0.858 3.022 0.986 ;
      RECT 2.976 0.922 3.086 0.986 ;
      RECT 2.938 0.922 3.086 0.944 ;
      RECT 2.63 0.835 2.976 0.925 ;
      RECT 3.03 0.17 3.12 0.345 ;
      RECT 2.32 0.17 2.41 0.345 ;
      RECT 2.32 0.17 3.12 0.26 ;
      RECT 1.84 0.205 1.93 1.135 ;
      RECT 1.84 0.669 2.01 0.809 ;
      RECT 0.78 1.14 1.416 1.23 ;
      RECT 0.78 1.14 1.462 1.207 ;
      RECT 1.378 1.121 1.508 1.161 ;
      RECT 0.78 0.43 0.87 1.23 ;
      RECT 1.416 1.079 1.508 1.161 ;
      RECT 1.462 1.033 1.554 1.115 ;
      RECT 1.508 0.987 1.6 1.069 ;
      RECT 1.508 0.987 1.646 1.023 ;
      RECT 1.554 0.941 1.65 0.998 ;
      RECT 1.6 0.895 1.696 0.973 ;
      RECT 1.646 0.87 1.65 0.998 ;
      RECT 1.65 0.765 1.74 0.928 ;
      RECT 0.78 0.43 0.92 0.52 ;
      RECT 1.275 0.823 1.365 1.018 ;
      RECT 1.24 0.423 1.33 0.862 ;
      RECT 1.225 0.635 1.33 0.837 ;
      RECT 1.275 0.383 1.386 0.446 ;
      RECT 1.33 0.346 1.34 0.474 ;
      RECT 1.34 0.205 1.43 0.401 ;
      RECT 1.321 0.355 1.43 0.401 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 1.02 0.935 1.16 1.05 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 1.02 0.17 1.11 1.05 ;
      RECT 1.02 0.405 1.15 0.545 ;
      RECT 0.045 0.445 0.64 0.535 ;
      RECT 0.55 0.17 0.64 0.535 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.55 0.17 1.11 0.26 ;
  END
END XNOR3X1H7R

MACRO XNOR3X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR3X1P4H7R 0 0 ;
  SIZE 4.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.2 1.48 ;
        RECT 3.29 1.05 3.38 1.48 ;
        RECT 2.81 1.035 2.9 1.48 ;
        RECT 1.575 1.2 1.665 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.2 0.08 ;
        RECT 3.76 -0.08 3.85 0.33 ;
        RECT 3.28 -0.08 3.37 0.345 ;
        RECT 1.59 -0.08 1.68 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.51 1.555 0.78 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.345 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.35 0.655 3.65 0.745 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.68 1.055 4.1 1.145 ;
        RECT 4.01 0.31 4.1 1.145 ;
      LAYER MET2 ;
        RECT 3.85 0.84 3.95 1.22 ;
      LAYER VIA1 ;
        RECT 3.855 1.055 3.945 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.335 0.435 2.425 1.015 ;
      RECT 3.214 0.855 3.92 0.945 ;
      RECT 3.83 0.595 3.92 0.945 ;
      RECT 3.201 0.81 3.214 0.939 ;
      RECT 3.155 0.781 3.201 0.909 ;
      RECT 3.109 0.735 3.155 0.863 ;
      RECT 3.109 0.836 3.252 0.863 ;
      RECT 3.063 0.689 3.109 0.817 ;
      RECT 3.017 0.643 3.063 0.771 ;
      RECT 2.979 0.689 3.109 0.729 ;
      RECT 2.335 0.62 3.017 0.71 ;
      RECT 2.07 0.435 2.665 0.525 ;
      RECT 2.525 0.35 2.665 0.525 ;
      RECT 2.07 0.205 2.16 0.525 ;
      RECT 2.775 0.44 3.6 0.53 ;
      RECT 3.51 0.205 3.6 0.53 ;
      RECT 2.775 0.35 2.915 0.53 ;
      RECT 2.07 1.105 2.72 1.195 ;
      RECT 2.63 0.835 2.72 1.195 ;
      RECT 3.04 0.967 3.13 1.135 ;
      RECT 2.07 1.035 2.16 1.195 ;
      RECT 3.022 0.89 3.04 1.018 ;
      RECT 2.976 0.858 3.022 0.986 ;
      RECT 2.976 0.922 3.086 0.986 ;
      RECT 2.938 0.922 3.086 0.944 ;
      RECT 2.63 0.835 2.976 0.925 ;
      RECT 3.03 0.17 3.12 0.345 ;
      RECT 2.32 0.17 2.41 0.345 ;
      RECT 2.32 0.17 3.12 0.26 ;
      RECT 1.84 0.205 1.93 1.135 ;
      RECT 1.84 0.669 2.01 0.809 ;
      RECT 0.78 1.14 1.416 1.23 ;
      RECT 0.78 1.14 1.462 1.207 ;
      RECT 1.378 1.121 1.508 1.161 ;
      RECT 0.78 0.43 0.87 1.23 ;
      RECT 1.416 1.079 1.508 1.161 ;
      RECT 1.462 1.033 1.554 1.115 ;
      RECT 1.508 0.987 1.6 1.069 ;
      RECT 1.508 0.987 1.646 1.023 ;
      RECT 1.554 0.941 1.65 0.998 ;
      RECT 1.6 0.895 1.696 0.973 ;
      RECT 1.646 0.87 1.65 0.998 ;
      RECT 1.65 0.765 1.74 0.928 ;
      RECT 0.78 0.43 0.92 0.52 ;
      RECT 1.275 0.823 1.365 1.018 ;
      RECT 1.24 0.418 1.33 0.862 ;
      RECT 1.225 0.635 1.33 0.837 ;
      RECT 1.275 0.378 1.386 0.441 ;
      RECT 1.33 0.341 1.34 0.469 ;
      RECT 1.34 0.205 1.43 0.396 ;
      RECT 1.321 0.35 1.43 0.396 ;
      RECT 0.045 1.01 0.185 1.1 ;
      RECT 1.02 0.935 1.16 1.05 ;
      RECT 0.045 0.23 0.135 1.1 ;
      RECT 1.02 0.17 1.11 1.05 ;
      RECT 1.02 0.405 1.15 0.545 ;
      RECT 0.045 0.44 0.64 0.53 ;
      RECT 0.55 0.17 0.64 0.53 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.55 0.17 1.11 0.26 ;
  END
END XNOR3X1P4H7R

MACRO XNOR3X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR3X2H7R 0 0 ;
  SIZE 4.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.6 1.48 ;
        RECT 3.96 1.235 4.1 1.48 ;
        RECT 3.29 1.05 3.38 1.48 ;
        RECT 2.81 1.035 2.9 1.48 ;
        RECT 1.575 1.2 1.665 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.6 0.08 ;
        RECT 4.26 -0.08 4.35 0.345 ;
        RECT 3.76 -0.08 3.85 0.33 ;
        RECT 3.28 -0.08 3.37 0.345 ;
        RECT 1.59 -0.08 1.68 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.505 1.555 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.345 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.35 0.655 3.65 0.745 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.68 1.055 4.1 1.145 ;
        RECT 4.01 0.22 4.1 1.145 ;
      LAYER MET2 ;
        RECT 3.85 0.84 3.95 1.22 ;
      LAYER VIA1 ;
        RECT 3.855 1.055 3.945 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.335 0.435 2.425 1.015 ;
      RECT 3.214 0.855 3.92 0.945 ;
      RECT 3.83 0.595 3.92 0.945 ;
      RECT 3.201 0.81 3.214 0.939 ;
      RECT 3.155 0.781 3.201 0.909 ;
      RECT 3.109 0.735 3.155 0.863 ;
      RECT 3.109 0.836 3.252 0.863 ;
      RECT 3.063 0.689 3.109 0.817 ;
      RECT 3.017 0.643 3.063 0.771 ;
      RECT 2.979 0.689 3.109 0.729 ;
      RECT 2.335 0.62 3.017 0.71 ;
      RECT 2.07 0.435 2.665 0.525 ;
      RECT 2.525 0.35 2.665 0.525 ;
      RECT 2.07 0.205 2.16 0.525 ;
      RECT 2.775 0.44 3.6 0.53 ;
      RECT 3.51 0.205 3.6 0.53 ;
      RECT 2.775 0.35 2.915 0.53 ;
      RECT 2.07 1.105 2.72 1.195 ;
      RECT 2.63 0.835 2.72 1.195 ;
      RECT 3.04 0.967 3.13 1.135 ;
      RECT 2.07 1.035 2.16 1.195 ;
      RECT 3.022 0.89 3.04 1.018 ;
      RECT 2.976 0.858 3.022 0.986 ;
      RECT 2.976 0.922 3.086 0.986 ;
      RECT 2.938 0.922 3.086 0.944 ;
      RECT 2.63 0.835 2.976 0.925 ;
      RECT 3.03 0.17 3.12 0.345 ;
      RECT 2.32 0.17 2.41 0.345 ;
      RECT 2.32 0.17 3.12 0.26 ;
      RECT 1.84 0.205 1.93 1.135 ;
      RECT 1.84 0.669 2.01 0.809 ;
      RECT 0.78 1.14 1.416 1.23 ;
      RECT 0.78 1.14 1.462 1.207 ;
      RECT 1.378 1.121 1.508 1.161 ;
      RECT 0.78 0.43 0.87 1.23 ;
      RECT 1.416 1.079 1.508 1.161 ;
      RECT 1.462 1.033 1.554 1.115 ;
      RECT 1.508 0.987 1.6 1.069 ;
      RECT 1.508 0.987 1.646 1.023 ;
      RECT 1.554 0.941 1.65 0.998 ;
      RECT 1.6 0.895 1.696 0.973 ;
      RECT 1.646 0.87 1.65 0.998 ;
      RECT 1.65 0.765 1.74 0.928 ;
      RECT 0.78 0.43 0.92 0.52 ;
      RECT 1.275 0.823 1.365 1.018 ;
      RECT 1.24 0.413 1.33 0.862 ;
      RECT 1.225 0.635 1.33 0.837 ;
      RECT 1.275 0.373 1.386 0.436 ;
      RECT 1.33 0.336 1.34 0.464 ;
      RECT 1.34 0.205 1.43 0.391 ;
      RECT 1.321 0.345 1.43 0.391 ;
      RECT 0.045 0.98 0.185 1.07 ;
      RECT 1.02 0.96 1.16 1.05 ;
      RECT 0.045 0.26 0.135 1.07 ;
      RECT 1.02 0.17 1.11 1.05 ;
      RECT 1.02 0.405 1.15 0.545 ;
      RECT 0.045 0.44 0.64 0.53 ;
      RECT 0.55 0.17 0.64 0.53 ;
      RECT 0.045 0.26 0.185 0.35 ;
      RECT 0.55 0.17 1.11 0.26 ;
  END
END XNOR3X2H7R

MACRO XNOR3X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR3X3H7R 0 0 ;
  SIZE 4.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.6 1.48 ;
        RECT 4.405 1.2 4.495 1.48 ;
        RECT 3.774 1.24 3.914 1.48 ;
        RECT 3.119 1.24 3.259 1.48 ;
        RECT 1.699 1.2 1.789 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.6 0.08 ;
        RECT 4.29 -0.08 4.38 0.33 ;
        RECT 3.679 -0.08 3.819 0.32 ;
        RECT 3.114 -0.08 3.204 0.33 ;
        RECT 1.59 -0.08 1.68 0.33 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.425 1.575 0.65 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.475 0.655 3.775 0.745 ;
      LAYER MET2 ;
        RECT 3.65 0.43 3.75 0.96 ;
      LAYER VIA1 ;
        RECT 3.655 0.655 3.745 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.115 1.05 4.33 1.14 ;
        RECT 4.24 0.507 4.33 1.14 ;
        RECT 4.191 0.462 4.286 0.541 ;
        RECT 4.132 0.437 4.24 0.466 ;
        RECT 4.237 0.507 4.33 0.566 ;
        RECT 4.132 0.413 4.237 0.466 ;
        RECT 4.086 0.367 4.191 0.436 ;
        RECT 4.145 0.462 4.286 0.495 ;
        RECT 4.04 0.225 4.145 0.39 ;
      LAYER MET2 ;
        RECT 4.05 0.18 4.15 0.56 ;
      LAYER VIA1 ;
        RECT 4.055 0.255 4.145 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.259 1.1 2.88 1.19 ;
      RECT 2.259 1.1 2.882 1.189 ;
      RECT 2.259 1.1 2.92 1.169 ;
      RECT 2.259 1.1 3.886 1.15 ;
      RECT 2.842 1.081 3.932 1.127 ;
      RECT 2.259 0.35 2.349 1.19 ;
      RECT 3.932 0.953 3.978 1.081 ;
      RECT 2.88 1.061 3.978 1.081 ;
      RECT 3.886 0.999 3.932 1.127 ;
      RECT 2.882 1.06 3.978 1.081 ;
      RECT 3.848 1.041 3.886 1.15 ;
      RECT 3.114 0.75 3.204 1.15 ;
      RECT 3.932 0.953 4.024 1.035 ;
      RECT 4.059 0.542 4.105 0.954 ;
      RECT 3.978 0.907 4.105 0.954 ;
      RECT 4.024 0.866 4.059 0.995 ;
      RECT 4.059 0.587 4.149 0.909 ;
      RECT 4.042 0.51 4.059 0.639 ;
      RECT 3.996 0.479 4.042 0.607 ;
      RECT 3.95 0.433 3.996 0.561 ;
      RECT 3.912 0.41 3.95 0.519 ;
      RECT 3.587 0.41 3.95 0.5 ;
      RECT 2.159 0.35 2.349 0.49 ;
      RECT 3.564 0.36 3.587 0.489 ;
      RECT 3.52 0.205 3.564 0.455 ;
      RECT 3.474 0.205 3.564 0.41 ;
      RECT 3.474 0.391 3.625 0.41 ;
      RECT 2.439 0.92 2.726 1.01 ;
      RECT 2.439 0.92 2.772 0.987 ;
      RECT 3.294 0.88 3.81 0.97 ;
      RECT 3.294 0.88 3.856 0.947 ;
      RECT 2.688 0.901 2.818 0.941 ;
      RECT 2.439 0.35 2.529 1.01 ;
      RECT 2.726 0.859 2.818 0.941 ;
      RECT 3.772 0.861 3.915 0.888 ;
      RECT 3.856 0.789 3.869 0.918 ;
      RECT 3.294 0.57 3.384 0.97 ;
      RECT 3.81 0.819 3.915 0.888 ;
      RECT 2.772 0.813 2.864 0.895 ;
      RECT 3.869 0.675 3.959 0.843 ;
      RECT 2.818 0.767 2.91 0.849 ;
      RECT 2.864 0.721 2.956 0.803 ;
      RECT 2.91 0.675 3.002 0.757 ;
      RECT 2.956 0.629 3.076 0.679 ;
      RECT 3.002 0.588 3.038 0.716 ;
      RECT 3.038 0.57 3.384 0.66 ;
      RECT 1.964 0.395 2.054 1.075 ;
      RECT 1.964 0.655 2.134 0.795 ;
      RECT 2.784 0.17 2.874 0.605 ;
      RECT 1.84 0.395 2.054 0.485 ;
      RECT 1.84 0.17 1.93 0.485 ;
      RECT 1.84 0.17 2.874 0.26 ;
      RECT 0.82 1.14 1.541 1.23 ;
      RECT 0.82 1.14 1.587 1.207 ;
      RECT 1.503 1.121 1.633 1.161 ;
      RECT 0.82 0.435 0.91 1.23 ;
      RECT 1.541 1.079 1.633 1.161 ;
      RECT 1.587 1.033 1.679 1.115 ;
      RECT 1.633 0.987 1.725 1.069 ;
      RECT 1.679 0.941 1.77 1.024 ;
      RECT 1.725 0.895 1.816 0.978 ;
      RECT 1.77 0.75 1.86 0.933 ;
      RECT 0.77 0.435 0.91 0.525 ;
      RECT 1.369 0.874 1.459 1.05 ;
      RECT 1.33 0.786 1.369 0.915 ;
      RECT 1.321 0.829 1.415 0.891 ;
      RECT 1.275 0.245 1.33 0.863 ;
      RECT 1.24 0.601 1.33 0.823 ;
      RECT 1.275 0.245 1.365 0.64 ;
      RECT 1.275 0.245 1.455 0.335 ;
      RECT 0.07 0.89 0.16 1.065 ;
      RECT 1.06 0.96 1.254 1.05 ;
      RECT 0.07 0.89 0.51 0.98 ;
      RECT 0.42 0.395 0.51 0.98 ;
      RECT 1.06 0.435 1.15 1.05 ;
      RECT 1.095 0.23 1.185 0.525 ;
      RECT 0.07 0.395 0.64 0.485 ;
      RECT 0.55 0.23 0.64 0.485 ;
      RECT 0.07 0.28 0.16 0.485 ;
      RECT 0.55 0.23 1.185 0.32 ;
  END
END XNOR3X3H7R

MACRO XNOR3X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR3X4H7R 0 0 ;
  SIZE 5 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5 1.48 ;
        RECT 4.59 1.035 4.68 1.48 ;
        RECT 3.974 1.225 4.114 1.48 ;
        RECT 3.399 1.225 3.539 1.48 ;
        RECT 1.979 1.2 2.069 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5 0.08 ;
        RECT 4.487 -0.08 4.577 0.33 ;
        RECT 3.984 -0.08 4.074 0.345 ;
        RECT 3.394 -0.08 3.484 0.33 ;
        RECT 1.909 -0.08 1.999 0.33 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.795 0.595 1.975 0.745 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.785 0.615 3.955 0.775 ;
      LAYER MET2 ;
        RECT 3.85 0.43 3.95 0.96 ;
      LAYER VIA1 ;
        RECT 3.855 0.655 3.945 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.405 0.455 4.827 0.545 ;
        RECT 4.737 0.255 4.827 0.545 ;
        RECT 4.315 1.06 4.495 1.15 ;
        RECT 4.405 0.455 4.495 1.15 ;
        RECT 4.37 0.439 4.482 0.489 ;
        RECT 4.324 0.401 4.451 0.448 ;
        RECT 4.28 0.36 4.405 0.403 ;
        RECT 4.28 0.32 4.37 0.403 ;
        RECT 4.234 0.19 4.324 0.358 ;
      LAYER MET2 ;
        RECT 4.45 0.225 4.55 0.76 ;
      LAYER VIA1 ;
        RECT 4.455 0.455 4.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.539 1.065 3.195 1.155 ;
      RECT 2.539 1.065 3.215 1.145 ;
      RECT 2.539 1.065 4.111 1.135 ;
      RECT 2.539 1.065 4.157 1.112 ;
      RECT 3.157 1.055 4.203 1.066 ;
      RECT 2.539 0.35 2.629 1.155 ;
      RECT 3.177 1.045 4.203 1.066 ;
      RECT 4.073 1.026 4.203 1.066 ;
      RECT 3.424 0.665 3.514 1.135 ;
      RECT 4.111 0.984 4.225 1.032 ;
      RECT 4.225 0.477 4.271 0.998 ;
      RECT 4.157 0.938 4.271 0.998 ;
      RECT 4.203 0.904 4.225 1.032 ;
      RECT 4.225 0.522 4.315 0.953 ;
      RECT 4.206 0.444 4.225 0.573 ;
      RECT 4.168 0.522 4.315 0.544 ;
      RECT 3.832 0.435 4.206 0.525 ;
      RECT 3.8 0.305 3.844 0.509 ;
      RECT 2.439 0.35 2.629 0.49 ;
      RECT 3.754 0.305 3.844 0.47 ;
      RECT 3.754 0.422 3.87 0.47 ;
      RECT 2.765 0.885 3.092 0.975 ;
      RECT 3.604 0.865 4.035 0.955 ;
      RECT 2.765 0.885 3.138 0.952 ;
      RECT 2.719 0.35 2.809 0.951 ;
      RECT 3.604 0.865 4.091 0.922 ;
      RECT 3.054 0.866 3.184 0.906 ;
      RECT 4.045 0.62 4.135 0.877 ;
      RECT 3.092 0.824 3.184 0.906 ;
      RECT 3.997 0.846 4.135 0.877 ;
      RECT 4.035 0.822 4.045 0.95 ;
      RECT 3.604 0.539 3.694 0.955 ;
      RECT 3.092 0.824 3.23 0.86 ;
      RECT 3.138 0.778 3.244 0.83 ;
      RECT 3.184 0.732 3.29 0.8 ;
      RECT 3.23 0.702 3.244 0.83 ;
      RECT 3.244 0.485 3.334 0.755 ;
      RECT 3.593 0.539 3.694 0.581 ;
      RECT 3.244 0.485 3.631 0.575 ;
      RECT 3.244 0.508 3.677 0.575 ;
      RECT 2.245 0.395 2.335 1.025 ;
      RECT 2.245 0.655 2.414 0.795 ;
      RECT 3.064 0.17 3.154 0.655 ;
      RECT 2.159 0.17 2.249 0.485 ;
      RECT 2.159 0.17 3.154 0.26 ;
      RECT 0.78 1.14 1.821 1.23 ;
      RECT 0.78 1.14 1.867 1.207 ;
      RECT 1.783 1.121 1.913 1.161 ;
      RECT 1.419 1.053 1.509 1.23 ;
      RECT 0.78 0.41 0.87 1.23 ;
      RECT 1.821 1.079 1.913 1.161 ;
      RECT 1.867 1.033 1.959 1.115 ;
      RECT 1.913 0.987 2.005 1.069 ;
      RECT 1.913 0.987 2.051 1.023 ;
      RECT 1.959 0.941 2.065 0.993 ;
      RECT 2.005 0.895 2.111 0.963 ;
      RECT 2.051 0.865 2.065 0.993 ;
      RECT 2.065 0.665 2.155 0.918 ;
      RECT 0.78 0.41 1.26 0.5 ;
      RECT 1.575 0.9 1.805 0.99 ;
      RECT 1.575 0.33 1.665 0.99 ;
      RECT 1.56 0.635 1.665 0.775 ;
      RECT 1.575 0.33 1.774 0.42 ;
      RECT 1.114 0.96 1.264 1.05 ;
      RECT 0.07 0.89 0.16 1.035 ;
      RECT 1.114 0.96 1.31 1.027 ;
      RECT 0.07 0.89 0.51 0.98 ;
      RECT 0.42 0.395 0.51 0.98 ;
      RECT 1.226 0.941 1.355 0.982 ;
      RECT 1.264 0.899 1.355 0.982 ;
      RECT 1.31 0.853 1.401 0.936 ;
      RECT 1.355 0.23 1.445 0.891 ;
      RECT 1.355 0.385 1.485 0.525 ;
      RECT 0.07 0.395 0.64 0.485 ;
      RECT 0.55 0.23 0.64 0.485 ;
      RECT 0.07 0.305 0.16 0.485 ;
      RECT 0.55 0.23 1.445 0.32 ;
  END
END XNOR3X4H7R

MACRO XNOR3X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR3X6H7R 0 0 ;
  SIZE 5.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5.2 1.48 ;
        RECT 4.605 1.2 4.695 1.48 ;
        RECT 3.974 1.225 4.114 1.48 ;
        RECT 3.399 1.225 3.539 1.48 ;
        RECT 1.979 1.2 2.069 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5.2 0.08 ;
        RECT 4.987 -0.08 5.077 0.345 ;
        RECT 4.487 -0.08 4.577 0.33 ;
        RECT 3.959 -0.08 4.099 0.32 ;
        RECT 3.394 -0.08 3.484 0.33 ;
        RECT 1.909 -0.08 1.999 0.33 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.8 0.595 1.95 0.775 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.784 0.605 3.945 0.775 ;
      LAYER MET2 ;
        RECT 3.85 0.43 3.95 0.96 ;
      LAYER VIA1 ;
        RECT 3.855 0.655 3.945 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.87 0.835 4.96 1.175 ;
        RECT 4.404 1.01 4.96 1.1 ;
        RECT 4.404 0.455 4.827 0.545 ;
        RECT 4.737 0.295 4.827 0.545 ;
        RECT 4.315 1.05 4.494 1.14 ;
        RECT 4.404 0.455 4.494 1.14 ;
        RECT 4.37 0.439 4.482 0.488 ;
        RECT 4.324 0.4 4.45 0.448 ;
        RECT 4.28 0.36 4.404 0.403 ;
        RECT 4.28 0.32 4.37 0.403 ;
        RECT 4.234 0.19 4.324 0.358 ;
      LAYER MET2 ;
        RECT 4.65 0.225 4.75 0.76 ;
      LAYER VIA1 ;
        RECT 4.655 0.455 4.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.539 1.065 3.195 1.155 ;
      RECT 2.539 1.065 3.215 1.145 ;
      RECT 2.539 1.065 4.101 1.135 ;
      RECT 2.539 1.065 4.147 1.112 ;
      RECT 3.157 1.055 4.193 1.066 ;
      RECT 2.539 0.35 2.629 1.155 ;
      RECT 3.177 1.045 4.193 1.066 ;
      RECT 4.063 1.026 4.193 1.066 ;
      RECT 3.424 0.665 3.514 1.135 ;
      RECT 4.101 0.984 4.224 1.028 ;
      RECT 4.224 0.477 4.27 0.989 ;
      RECT 4.147 0.938 4.27 0.989 ;
      RECT 4.193 0.899 4.224 1.028 ;
      RECT 4.224 0.522 4.314 0.944 ;
      RECT 4.195 0.439 4.224 0.568 ;
      RECT 4.157 0.425 4.195 0.534 ;
      RECT 3.882 0.425 4.195 0.515 ;
      RECT 3.844 0.368 3.882 0.496 ;
      RECT 2.439 0.35 2.629 0.49 ;
      RECT 3.8 0.406 3.92 0.455 ;
      RECT 3.754 0.205 3.844 0.41 ;
      RECT 2.719 0.885 3.092 0.975 ;
      RECT 3.604 0.865 4.025 0.955 ;
      RECT 2.719 0.885 3.138 0.952 ;
      RECT 3.604 0.865 4.09 0.913 ;
      RECT 3.054 0.866 3.184 0.906 ;
      RECT 2.719 0.35 2.809 0.975 ;
      RECT 4.044 0.62 4.134 0.868 ;
      RECT 3.092 0.824 3.184 0.906 ;
      RECT 3.987 0.846 4.134 0.868 ;
      RECT 4.025 0.817 4.044 0.946 ;
      RECT 3.604 0.539 3.694 0.955 ;
      RECT 3.092 0.824 3.23 0.86 ;
      RECT 3.138 0.778 3.244 0.83 ;
      RECT 3.184 0.732 3.29 0.8 ;
      RECT 3.23 0.702 3.244 0.83 ;
      RECT 3.244 0.485 3.334 0.755 ;
      RECT 3.593 0.539 3.694 0.581 ;
      RECT 3.244 0.485 3.631 0.575 ;
      RECT 3.244 0.508 3.677 0.575 ;
      RECT 2.244 0.395 2.334 1.015 ;
      RECT 2.244 0.655 2.414 0.795 ;
      RECT 3.064 0.17 3.154 0.655 ;
      RECT 2.159 0.17 2.249 0.485 ;
      RECT 2.159 0.17 3.154 0.26 ;
      RECT 0.78 1.14 1.821 1.23 ;
      RECT 0.78 1.14 1.867 1.207 ;
      RECT 1.783 1.121 1.913 1.161 ;
      RECT 1.419 1.028 1.509 1.23 ;
      RECT 0.78 0.41 0.87 1.23 ;
      RECT 1.821 1.079 1.913 1.161 ;
      RECT 1.867 1.033 1.959 1.115 ;
      RECT 1.913 0.987 2.005 1.069 ;
      RECT 1.913 0.987 2.051 1.023 ;
      RECT 1.959 0.941 2.064 0.994 ;
      RECT 2.005 0.895 2.11 0.964 ;
      RECT 2.051 0.865 2.064 0.994 ;
      RECT 2.064 0.69 2.154 0.919 ;
      RECT 0.78 0.41 1.26 0.5 ;
      RECT 1.62 0.9 1.805 0.99 ;
      RECT 1.62 0.33 1.71 0.99 ;
      RECT 1.535 0.66 1.71 0.75 ;
      RECT 1.62 0.33 1.774 0.42 ;
      RECT 1.114 0.96 1.264 1.05 ;
      RECT 0.07 0.89 0.16 1.035 ;
      RECT 1.114 0.96 1.31 1.027 ;
      RECT 0.07 0.89 0.51 0.98 ;
      RECT 0.42 0.395 0.51 0.98 ;
      RECT 1.226 0.941 1.355 0.982 ;
      RECT 1.264 0.899 1.355 0.982 ;
      RECT 1.31 0.853 1.401 0.936 ;
      RECT 1.355 0.23 1.445 0.891 ;
      RECT 1.355 0.385 1.485 0.525 ;
      RECT 0.07 0.395 0.64 0.485 ;
      RECT 0.55 0.23 0.64 0.485 ;
      RECT 0.07 0.305 0.16 0.485 ;
      RECT 0.55 0.23 1.445 0.32 ;
  END
END XNOR3X6H7R

MACRO XOR2X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2X0P5H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.575 1.2 1.665 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.59 -0.08 1.68 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.505 1.555 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.765 0.375 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.84 0.205 1.945 0.375 ;
        RECT 1.84 0.205 1.93 1.135 ;
      LAYER MET2 ;
        RECT 1.85 0.18 1.95 0.56 ;
      LAYER VIA1 ;
        RECT 1.855 0.255 1.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.78 1.14 1.415 1.23 ;
      RECT 0.78 1.14 1.461 1.207 ;
      RECT 1.377 1.121 1.507 1.161 ;
      RECT 0.78 0.43 0.87 1.23 ;
      RECT 1.415 1.079 1.507 1.161 ;
      RECT 1.461 1.033 1.553 1.115 ;
      RECT 1.507 0.987 1.599 1.069 ;
      RECT 1.507 0.987 1.645 1.023 ;
      RECT 1.553 0.941 1.65 0.998 ;
      RECT 1.599 0.895 1.696 0.972 ;
      RECT 1.645 0.869 1.65 0.998 ;
      RECT 1.65 0.765 1.74 0.927 ;
      RECT 0.78 0.43 0.92 0.52 ;
      RECT 1.275 0.823 1.365 1.018 ;
      RECT 1.24 0.393 1.33 0.862 ;
      RECT 1.23 0.635 1.33 0.839 ;
      RECT 1.275 0.353 1.386 0.416 ;
      RECT 1.33 0.316 1.34 0.444 ;
      RECT 1.34 0.205 1.43 0.371 ;
      RECT 1.321 0.325 1.43 0.371 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 1.02 0.96 1.16 1.05 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 1.02 0.25 1.11 1.05 ;
      RECT 1.02 0.405 1.15 0.545 ;
      RECT 0.045 0.445 0.64 0.535 ;
      RECT 0.55 0.25 0.64 0.535 ;
      RECT 0.55 0.25 1.11 0.34 ;
      RECT 0.045 0.23 0.185 0.32 ;
  END
END XOR2X0P5H7R

MACRO XOR2X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2X0P7H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.575 1.2 1.665 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.59 -0.08 1.68 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.475 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.345 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.84 0.225 1.945 0.375 ;
        RECT 1.84 0.225 1.93 1.103 ;
      LAYER MET2 ;
        RECT 1.85 0.18 1.95 0.56 ;
      LAYER VIA1 ;
        RECT 1.855 0.255 1.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.78 1.14 1.416 1.23 ;
      RECT 0.78 1.14 1.462 1.207 ;
      RECT 1.378 1.121 1.508 1.161 ;
      RECT 0.78 0.43 0.87 1.23 ;
      RECT 1.416 1.079 1.508 1.161 ;
      RECT 1.462 1.033 1.554 1.115 ;
      RECT 1.508 0.987 1.6 1.069 ;
      RECT 1.508 0.987 1.646 1.023 ;
      RECT 1.554 0.941 1.66 0.993 ;
      RECT 1.6 0.895 1.706 0.963 ;
      RECT 1.646 0.865 1.66 0.993 ;
      RECT 1.66 0.753 1.75 0.918 ;
      RECT 0.78 0.43 0.92 0.52 ;
      RECT 1.275 0.823 1.365 1.018 ;
      RECT 1.241 0.388 1.33 0.862 ;
      RECT 1.24 0.405 1.33 0.845 ;
      RECT 1.225 0.635 1.33 0.837 ;
      RECT 1.33 0.311 1.34 0.439 ;
      RECT 1.275 0.348 1.386 0.411 ;
      RECT 1.321 0.32 1.33 1.018 ;
      RECT 1.34 0.205 1.429 0.367 ;
      RECT 1.34 0.205 1.43 0.345 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 1.02 0.96 1.16 1.05 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 1.02 0.17 1.11 1.05 ;
      RECT 1.02 0.405 1.15 0.545 ;
      RECT 0.045 0.445 0.64 0.535 ;
      RECT 0.55 0.17 0.64 0.535 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.55 0.17 1.11 0.26 ;
  END
END XOR2X0P7H7R

MACRO XOR2X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2X1H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.575 1.2 1.665 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.59 -0.08 1.68 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.475 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.345 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.815 0.96 1.955 1.05 ;
        RECT 1.855 0.29 1.955 1.05 ;
        RECT 1.815 0.29 1.955 0.38 ;
      LAYER MET2 ;
        RECT 1.85 0.625 1.95 1.16 ;
      LAYER VIA1 ;
        RECT 1.855 0.855 1.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.78 1.14 1.414 1.23 ;
      RECT 0.78 1.14 1.46 1.207 ;
      RECT 1.376 1.121 1.506 1.161 ;
      RECT 0.78 0.43 0.87 1.23 ;
      RECT 1.414 1.079 1.506 1.161 ;
      RECT 1.46 1.033 1.552 1.115 ;
      RECT 1.506 0.987 1.598 1.069 ;
      RECT 1.552 0.941 1.644 1.023 ;
      RECT 1.598 0.895 1.721 0.946 ;
      RECT 1.644 0.856 1.675 0.985 ;
      RECT 1.675 0.705 1.765 0.901 ;
      RECT 0.78 0.43 0.92 0.52 ;
      RECT 1.275 0.823 1.365 1.018 ;
      RECT 1.241 0.388 1.33 0.862 ;
      RECT 1.24 0.405 1.33 0.845 ;
      RECT 1.225 0.635 1.33 0.837 ;
      RECT 1.33 0.311 1.34 0.439 ;
      RECT 1.275 0.348 1.386 0.411 ;
      RECT 1.321 0.32 1.33 1.018 ;
      RECT 1.34 0.205 1.429 0.367 ;
      RECT 1.34 0.205 1.43 0.345 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 1.02 0.935 1.16 1.05 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 1.02 0.17 1.11 1.05 ;
      RECT 1.02 0.405 1.15 0.545 ;
      RECT 0.045 0.445 0.64 0.535 ;
      RECT 0.55 0.17 0.64 0.535 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.55 0.17 1.11 0.26 ;
  END
END XOR2X1H7R

MACRO XOR2X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2X1P4H7R 0 0 ;
  SIZE 2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2 1.48 ;
        RECT 1.575 1.2 1.665 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2 0.08 ;
        RECT 1.59 -0.08 1.68 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.445 0.505 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.345 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.815 0.96 1.955 1.05 ;
        RECT 1.855 0.326 1.955 1.05 ;
        RECT 1.815 0.326 1.955 0.416 ;
      LAYER MET2 ;
        RECT 1.85 0.625 1.95 1.16 ;
      LAYER VIA1 ;
        RECT 1.855 0.855 1.945 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.78 1.14 1.414 1.23 ;
      RECT 0.78 1.14 1.46 1.207 ;
      RECT 1.376 1.121 1.506 1.161 ;
      RECT 0.78 0.43 0.87 1.23 ;
      RECT 1.414 1.079 1.506 1.161 ;
      RECT 1.46 1.033 1.552 1.115 ;
      RECT 1.506 0.987 1.598 1.069 ;
      RECT 1.552 0.941 1.644 1.023 ;
      RECT 1.598 0.895 1.721 0.946 ;
      RECT 1.644 0.856 1.675 0.985 ;
      RECT 1.675 0.661 1.765 0.901 ;
      RECT 0.78 0.43 0.92 0.52 ;
      RECT 1.275 0.823 1.365 1.018 ;
      RECT 1.24 0.418 1.33 0.862 ;
      RECT 1.215 0.635 1.33 0.832 ;
      RECT 1.275 0.378 1.386 0.441 ;
      RECT 1.33 0.341 1.34 0.469 ;
      RECT 1.34 0.205 1.43 0.396 ;
      RECT 1.321 0.35 1.43 0.396 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 1.02 0.96 1.16 1.05 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 1.02 0.17 1.11 1.05 ;
      RECT 1.02 0.405 1.15 0.545 ;
      RECT 0.045 0.445 0.64 0.535 ;
      RECT 0.55 0.17 0.64 0.535 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.55 0.17 1.11 0.26 ;
  END
END XOR2X1P4H7R

MACRO XOR2X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2X2H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 2.09 1.035 2.18 1.48 ;
        RECT 1.575 1.2 1.665 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 2.09 -0.08 2.18 0.345 ;
        RECT 1.59 -0.08 1.68 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.48 1.545 0.78 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.625 0.345 0.85 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.84 0.22 1.945 1.12 ;
      LAYER MET2 ;
        RECT 1.85 0.18 1.95 0.56 ;
      LAYER VIA1 ;
        RECT 1.855 0.255 1.945 0.345 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.78 1.14 1.414 1.23 ;
      RECT 0.78 1.14 1.46 1.207 ;
      RECT 1.376 1.121 1.506 1.161 ;
      RECT 0.78 0.43 0.92 1.23 ;
      RECT 1.414 1.079 1.506 1.161 ;
      RECT 1.46 1.033 1.552 1.115 ;
      RECT 1.506 0.987 1.598 1.069 ;
      RECT 1.506 0.987 1.644 1.023 ;
      RECT 1.552 0.941 1.65 0.997 ;
      RECT 1.598 0.895 1.696 0.971 ;
      RECT 1.644 0.869 1.65 0.997 ;
      RECT 1.65 0.76 1.74 0.926 ;
      RECT 1.275 0.823 1.365 1.018 ;
      RECT 1.24 0.403 1.33 0.862 ;
      RECT 1.225 0.635 1.33 0.837 ;
      RECT 1.275 0.363 1.386 0.426 ;
      RECT 1.33 0.326 1.34 0.454 ;
      RECT 1.34 0.205 1.43 0.381 ;
      RECT 1.321 0.335 1.43 0.381 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 1.02 0.96 1.16 1.05 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 1.02 0.17 1.11 1.05 ;
      RECT 1.02 0.405 1.15 0.545 ;
      RECT 0.045 0.445 0.64 0.535 ;
      RECT 0.55 0.17 0.64 0.535 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.55 0.17 1.11 0.26 ;
  END
END XOR2X2H7R

MACRO XOR2X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2X3H7R 0 0 ;
  SIZE 2.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.4 1.48 ;
        RECT 2.105 1.035 2.195 1.48 ;
        RECT 1.59 1.2 1.68 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.4 0.08 ;
        RECT 2.09 -0.08 2.18 0.345 ;
        RECT 1.575 -0.08 1.665 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.445 0.55 1.565 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.24 0.715 0.345 0.975 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.855 0.855 2.145 0.945 ;
        RECT 2.055 0.435 2.145 0.945 ;
        RECT 1.84 0.435 2.145 0.525 ;
        RECT 1.855 0.855 1.945 1.025 ;
        RECT 1.84 0.295 1.93 0.525 ;
      LAYER MET2 ;
        RECT 2.05 0.43 2.15 0.96 ;
      LAYER VIA1 ;
        RECT 2.055 0.655 2.145 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.78 1.14 1.429 1.23 ;
      RECT 0.78 1.14 1.475 1.207 ;
      RECT 1.391 1.121 1.521 1.161 ;
      RECT 0.78 0.43 0.87 1.23 ;
      RECT 1.429 1.079 1.521 1.161 ;
      RECT 1.475 1.033 1.567 1.115 ;
      RECT 1.521 0.987 1.613 1.069 ;
      RECT 1.521 0.987 1.659 1.023 ;
      RECT 1.567 0.941 1.675 0.992 ;
      RECT 1.613 0.895 1.721 0.961 ;
      RECT 1.659 0.864 1.675 0.992 ;
      RECT 1.675 0.675 1.765 0.916 ;
      RECT 1.675 0.675 1.885 0.765 ;
      RECT 0.78 0.43 0.92 0.52 ;
      RECT 1.29 0.839 1.38 1.018 ;
      RECT 1.286 0.348 1.33 0.877 ;
      RECT 1.24 0.373 1.33 0.852 ;
      RECT 1.24 0.814 1.376 0.852 ;
      RECT 1.325 0.205 1.376 0.411 ;
      RECT 1.325 0.205 1.415 0.369 ;
      RECT 1.29 0.328 1.415 0.369 ;
      RECT 0.045 1.05 0.185 1.14 ;
      RECT 1.035 0.96 1.175 1.05 ;
      RECT 0.045 0.23 0.135 1.14 ;
      RECT 1.035 0.17 1.15 1.05 ;
      RECT 0.045 0.5 0.64 0.59 ;
      RECT 0.55 0.17 0.64 0.59 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.55 0.17 1.15 0.26 ;
  END
END XOR2X3H7R

MACRO XOR2X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2X4H7R 0 0 ;
  SIZE 2.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 2.6 1.48 ;
        RECT 2.221 1.055 2.311 1.48 ;
        RECT 1.656 1.2 1.746 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 2.6 0.08 ;
        RECT 2.066 -0.08 2.206 0.305 ;
        RECT 1.591 -0.08 1.681 0.33 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.425 1.59 0.625 ;
      LAYER MET2 ;
        RECT 1.45 0.23 1.55 0.76 ;
      LAYER VIA1 ;
        RECT 1.455 0.455 1.545 0.545 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.841 0.395 2.431 0.485 ;
        RECT 2.341 0.255 2.431 0.485 ;
        RECT 1.946 0.835 2.345 0.925 ;
        RECT 2.255 0.395 2.345 0.925 ;
        RECT 1.841 0.27 1.931 0.485 ;
      LAYER MET2 ;
        RECT 2.25 0.43 2.35 0.96 ;
      LAYER VIA1 ;
        RECT 2.255 0.655 2.345 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.82 1.14 1.479 1.23 ;
      RECT 0.82 1.14 1.525 1.207 ;
      RECT 1.441 1.121 1.571 1.161 ;
      RECT 0.82 0.43 0.91 1.23 ;
      RECT 1.479 1.079 1.571 1.161 ;
      RECT 1.525 1.033 1.617 1.115 ;
      RECT 1.571 0.987 1.663 1.069 ;
      RECT 1.617 0.941 1.709 1.023 ;
      RECT 1.663 0.895 1.786 0.946 ;
      RECT 1.709 0.856 1.74 0.985 ;
      RECT 1.74 0.605 1.83 0.901 ;
      RECT 1.74 0.605 2.086 0.695 ;
      RECT 0.82 0.43 0.96 0.52 ;
      RECT 1.326 0.835 1.416 1.018 ;
      RECT 1.321 0.835 1.416 0.889 ;
      RECT 1.275 0.795 1.381 0.863 ;
      RECT 1.245 0.62 1.335 0.825 ;
      RECT 1.275 0.23 1.365 0.658 ;
      RECT 1.275 0.23 1.456 0.32 ;
      RECT 1.065 0.96 1.211 1.05 ;
      RECT 0.07 0.89 0.16 1.035 ;
      RECT 0.07 0.89 0.51 0.98 ;
      RECT 0.42 0.395 0.51 0.98 ;
      RECT 1.065 0.25 1.155 1.05 ;
      RECT 1.065 0.25 1.185 0.545 ;
      RECT 0.07 0.395 0.64 0.485 ;
      RECT 0.55 0.25 0.64 0.485 ;
      RECT 0.07 0.305 0.16 0.485 ;
      RECT 0.55 0.25 1.185 0.34 ;
  END
END XOR2X4H7R

MACRO XOR2X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2X6H7R 0 0 ;
  SIZE 3 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 3 1.48 ;
        RECT 2.514 1.07 2.604 1.48 ;
        RECT 1.949 1.2 2.039 1.48 ;
        RECT 0.57 1.07 0.66 1.48 ;
        RECT 0.07 1.055 0.16 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 3 0.08 ;
        RECT 2.825 -0.08 2.915 0.345 ;
        RECT 2.3 -0.08 2.44 0.305 ;
        RECT 1.825 -0.08 1.915 0.33 ;
        RECT 0.545 -0.08 0.685 0.305 ;
        RECT 0.07 -0.08 0.16 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.745 0.625 1.945 0.775 ;
      LAYER MET2 ;
        RECT 1.85 0.425 1.95 0.96 ;
      LAYER VIA1 ;
        RECT 1.855 0.655 1.945 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.195 0.655 0.535 0.745 ;
      LAYER MET2 ;
        RECT 0.25 0.425 0.35 0.96 ;
      LAYER VIA1 ;
        RECT 0.255 0.655 0.345 0.745 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.239 0.855 2.879 0.945 ;
        RECT 2.575 0.22 2.665 0.945 ;
        RECT 2.075 0.395 2.665 0.485 ;
        RECT 2.075 0.32 2.165 0.485 ;
      LAYER MET2 ;
        RECT 2.65 0.63 2.75 1.16 ;
      LAYER VIA1 ;
        RECT 2.655 0.855 2.745 0.945 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.07 1.14 1.791 1.23 ;
      RECT 1.07 1.14 1.837 1.207 ;
      RECT 1.753 1.121 1.873 1.166 ;
      RECT 1.07 0.43 1.16 1.23 ;
      RECT 1.791 1.079 1.911 1.129 ;
      RECT 1.837 1.038 1.873 1.166 ;
      RECT 2.035 0.62 2.125 1.11 ;
      RECT 1.873 1.02 2.125 1.11 ;
      RECT 2.035 0.62 2.375 0.71 ;
      RECT 1.07 0.43 1.21 0.52 ;
      RECT 1.619 0.874 1.709 1.05 ;
      RECT 1.58 0.786 1.619 0.915 ;
      RECT 1.571 0.829 1.665 0.891 ;
      RECT 1.525 0.23 1.58 0.863 ;
      RECT 1.49 0.616 1.58 0.823 ;
      RECT 1.525 0.23 1.615 0.655 ;
      RECT 1.525 0.23 1.69 0.32 ;
      RECT 0.32 0.89 0.41 1.14 ;
      RECT 1.3 0.96 1.504 1.05 ;
      RECT 0.32 0.89 0.76 0.98 ;
      RECT 0.67 0.395 0.76 0.98 ;
      RECT 1.3 0.455 1.39 1.05 ;
      RECT 1.345 0.25 1.435 0.545 ;
      RECT 0.32 0.395 0.89 0.485 ;
      RECT 0.8 0.25 0.89 0.485 ;
      RECT 0.32 0.22 0.41 0.485 ;
      RECT 0.8 0.25 1.435 0.34 ;
  END
END XOR2X6H7R

MACRO XOR3X0P5H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR3X0P5H7R 0 0 ;
  SIZE 4.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.2 1.48 ;
        RECT 3.29 1.05 3.38 1.48 ;
        RECT 2.81 1.035 2.9 1.48 ;
        RECT 1.575 1.2 1.665 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.2 0.08 ;
        RECT 3.76 -0.08 3.85 0.33 ;
        RECT 3.28 -0.08 3.37 0.345 ;
        RECT 1.59 -0.08 1.68 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.505 1.555 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.765 0.375 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.225 0.81 3.425 0.945 ;
      LAYER MET2 ;
        RECT 3.25 0.63 3.35 1.16 ;
      LAYER VIA1 ;
        RECT 3.255 0.855 3.345 0.945 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.68 1.055 4.1 1.145 ;
        RECT 4.01 0.205 4.1 1.145 ;
      LAYER MET2 ;
        RECT 3.85 0.84 3.95 1.22 ;
      LAYER VIA1 ;
        RECT 3.855 1.055 3.945 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.335 0.435 2.425 1.05 ;
      RECT 3.83 0.62 3.92 0.76 ;
      RECT 2.335 0.62 3.92 0.71 ;
      RECT 2.07 0.435 2.665 0.525 ;
      RECT 2.525 0.35 2.665 0.525 ;
      RECT 2.07 0.205 2.16 0.525 ;
      RECT 2.775 0.44 3.6 0.53 ;
      RECT 3.51 0.205 3.6 0.53 ;
      RECT 2.775 0.35 2.915 0.53 ;
      RECT 2.07 1.14 2.72 1.23 ;
      RECT 2.63 0.835 2.72 1.23 ;
      RECT 2.07 1.035 2.16 1.23 ;
      RECT 3.04 0.835 3.13 1.135 ;
      RECT 2.63 0.835 3.13 0.925 ;
      RECT 3.03 0.17 3.12 0.345 ;
      RECT 2.32 0.17 2.41 0.345 ;
      RECT 2.32 0.17 3.12 0.26 ;
      RECT 1.84 0.205 1.93 1.135 ;
      RECT 1.84 0.694 2.105 0.784 ;
      RECT 0.78 1.14 1.416 1.23 ;
      RECT 0.78 1.14 1.462 1.207 ;
      RECT 1.378 1.121 1.508 1.161 ;
      RECT 0.78 0.35 0.87 1.23 ;
      RECT 1.416 1.079 1.508 1.161 ;
      RECT 1.462 1.033 1.554 1.115 ;
      RECT 1.508 0.987 1.6 1.069 ;
      RECT 1.508 0.987 1.646 1.023 ;
      RECT 1.554 0.941 1.65 0.998 ;
      RECT 1.6 0.895 1.696 0.973 ;
      RECT 1.646 0.87 1.65 0.998 ;
      RECT 1.65 0.765 1.74 0.928 ;
      RECT 0.78 0.35 0.925 0.44 ;
      RECT 1.275 0.712 1.365 1.018 ;
      RECT 1.241 0.672 1.331 0.75 ;
      RECT 1.195 0.452 1.285 0.71 ;
      RECT 1.195 0.452 1.331 0.49 ;
      RECT 1.241 0.412 1.34 0.463 ;
      RECT 1.275 0.39 1.386 0.435 ;
      RECT 1.331 0.334 1.34 0.463 ;
      RECT 1.34 0.205 1.43 0.39 ;
      RECT 1.285 0.362 1.43 0.39 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 1.015 0.84 1.16 0.93 ;
      RECT 1.015 0.17 1.105 0.93 ;
      RECT 0.045 0.445 0.64 0.535 ;
      RECT 0.55 0.17 0.64 0.535 ;
      RECT 1.015 0.17 1.18 0.345 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.55 0.17 1.18 0.26 ;
  END
END XOR3X0P5H7R

MACRO XOR3X0P7H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR3X0P7H7R 0 0 ;
  SIZE 4.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.2 1.48 ;
        RECT 3.29 1.05 3.38 1.48 ;
        RECT 2.81 1.035 2.9 1.48 ;
        RECT 1.575 1.2 1.665 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.2 0.08 ;
        RECT 3.76 -0.08 3.85 0.33 ;
        RECT 3.28 -0.08 3.37 0.345 ;
        RECT 1.59 -0.08 1.68 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.475 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.765 0.375 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.225 0.8 3.415 0.945 ;
      LAYER MET2 ;
        RECT 3.25 0.63 3.35 1.16 ;
      LAYER VIA1 ;
        RECT 3.255 0.855 3.345 0.945 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.68 1.055 4.1 1.145 ;
        RECT 4.01 0.229 4.1 1.145 ;
      LAYER MET2 ;
        RECT 3.85 0.84 3.95 1.22 ;
      LAYER VIA1 ;
        RECT 3.855 1.055 3.945 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.335 0.435 2.43 1.015 ;
      RECT 3.83 0.62 3.92 0.76 ;
      RECT 2.335 0.62 3.92 0.71 ;
      RECT 2.07 0.435 2.665 0.525 ;
      RECT 2.525 0.35 2.665 0.525 ;
      RECT 2.07 0.205 2.16 0.525 ;
      RECT 2.775 0.44 3.6 0.53 ;
      RECT 3.51 0.205 3.6 0.53 ;
      RECT 2.775 0.35 2.915 0.53 ;
      RECT 2.07 1.14 2.72 1.23 ;
      RECT 2.63 0.835 2.72 1.23 ;
      RECT 2.07 1.035 2.16 1.23 ;
      RECT 3.04 0.835 3.13 1.135 ;
      RECT 2.63 0.835 3.13 0.925 ;
      RECT 3.03 0.17 3.12 0.345 ;
      RECT 2.32 0.17 2.41 0.345 ;
      RECT 2.32 0.17 3.12 0.26 ;
      RECT 1.84 0.205 1.93 1.135 ;
      RECT 1.84 0.685 2.035 0.775 ;
      RECT 0.78 1.11 1.446 1.2 ;
      RECT 0.78 1.11 1.492 1.177 ;
      RECT 1.408 1.091 1.538 1.131 ;
      RECT 0.78 0.35 0.87 1.2 ;
      RECT 1.446 1.049 1.538 1.131 ;
      RECT 1.492 1.003 1.584 1.085 ;
      RECT 1.492 1.003 1.63 1.039 ;
      RECT 1.538 0.957 1.65 1.006 ;
      RECT 1.584 0.911 1.696 0.973 ;
      RECT 1.63 0.878 1.65 1.006 ;
      RECT 1.65 0.765 1.74 0.928 ;
      RECT 0.78 0.35 0.925 0.44 ;
      RECT 1.275 0.712 1.365 1.018 ;
      RECT 1.241 0.672 1.331 0.75 ;
      RECT 1.195 0.437 1.285 0.71 ;
      RECT 1.195 0.437 1.331 0.475 ;
      RECT 1.241 0.397 1.34 0.448 ;
      RECT 1.275 0.375 1.386 0.42 ;
      RECT 1.331 0.319 1.34 0.448 ;
      RECT 1.34 0.205 1.43 0.375 ;
      RECT 1.285 0.347 1.43 0.375 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 1.015 0.865 1.16 0.955 ;
      RECT 1.015 0.17 1.105 0.955 ;
      RECT 0.045 0.445 0.64 0.535 ;
      RECT 0.55 0.17 0.64 0.535 ;
      RECT 1.015 0.17 1.18 0.345 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.55 0.17 1.18 0.26 ;
  END
END XOR3X0P7H7R

MACRO XOR3X1H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR3X1H7R 0 0 ;
  SIZE 4.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.2 1.48 ;
        RECT 3.29 1.05 3.38 1.48 ;
        RECT 2.81 1.035 2.9 1.48 ;
        RECT 1.575 1.2 1.665 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.2 0.08 ;
        RECT 3.76 -0.08 3.85 0.33 ;
        RECT 3.28 -0.08 3.37 0.345 ;
        RECT 1.59 -0.08 1.68 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.475 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.765 0.375 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.35 0.655 3.65 0.745 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.68 1.055 4.1 1.145 ;
        RECT 4.01 0.265 4.1 1.145 ;
      LAYER MET2 ;
        RECT 3.85 0.84 3.95 1.22 ;
      LAYER VIA1 ;
        RECT 3.855 1.055 3.945 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.335 0.435 2.425 1.015 ;
      RECT 3.194 0.835 3.92 0.925 ;
      RECT 3.83 0.705 3.92 0.925 ;
      RECT 3.155 0.777 3.194 0.906 ;
      RECT 3.109 0.735 3.155 0.863 ;
      RECT 3.109 0.816 3.232 0.863 ;
      RECT 3.063 0.689 3.109 0.817 ;
      RECT 3.017 0.643 3.063 0.771 ;
      RECT 2.979 0.689 3.109 0.729 ;
      RECT 2.335 0.62 3.017 0.71 ;
      RECT 2.07 0.435 2.665 0.525 ;
      RECT 2.525 0.35 2.665 0.525 ;
      RECT 2.07 0.205 2.16 0.525 ;
      RECT 2.775 0.44 3.6 0.53 ;
      RECT 3.51 0.205 3.6 0.53 ;
      RECT 2.775 0.35 2.915 0.53 ;
      RECT 2.07 1.105 2.72 1.195 ;
      RECT 2.63 0.835 2.72 1.195 ;
      RECT 3.04 0.967 3.13 1.135 ;
      RECT 2.07 1.035 2.16 1.195 ;
      RECT 3.022 0.89 3.04 1.018 ;
      RECT 2.976 0.858 3.022 0.986 ;
      RECT 2.976 0.922 3.086 0.986 ;
      RECT 2.938 0.922 3.086 0.944 ;
      RECT 2.63 0.835 2.976 0.925 ;
      RECT 3.03 0.17 3.12 0.345 ;
      RECT 2.32 0.17 2.41 0.345 ;
      RECT 2.32 0.17 3.12 0.26 ;
      RECT 1.84 0.205 1.93 1.135 ;
      RECT 1.84 0.694 2.035 0.784 ;
      RECT 0.78 1.14 1.416 1.23 ;
      RECT 0.78 1.14 1.462 1.207 ;
      RECT 1.378 1.121 1.508 1.161 ;
      RECT 0.78 0.35 0.87 1.23 ;
      RECT 1.416 1.079 1.508 1.161 ;
      RECT 1.462 1.033 1.554 1.115 ;
      RECT 1.508 0.987 1.6 1.069 ;
      RECT 1.508 0.987 1.646 1.023 ;
      RECT 1.554 0.941 1.65 0.998 ;
      RECT 1.6 0.895 1.696 0.973 ;
      RECT 1.646 0.87 1.65 0.998 ;
      RECT 1.65 0.765 1.74 0.928 ;
      RECT 0.78 0.35 0.925 0.44 ;
      RECT 1.275 0.712 1.365 1.018 ;
      RECT 1.241 0.672 1.331 0.75 ;
      RECT 1.195 0.437 1.285 0.71 ;
      RECT 1.195 0.437 1.331 0.475 ;
      RECT 1.241 0.397 1.34 0.448 ;
      RECT 1.275 0.375 1.386 0.42 ;
      RECT 1.331 0.319 1.34 0.448 ;
      RECT 1.34 0.205 1.43 0.375 ;
      RECT 1.285 0.347 1.43 0.375 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 1.015 0.84 1.16 0.93 ;
      RECT 1.015 0.17 1.105 0.93 ;
      RECT 0.045 0.445 0.64 0.535 ;
      RECT 0.55 0.17 0.64 0.535 ;
      RECT 1.015 0.17 1.18 0.345 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.55 0.17 1.18 0.26 ;
  END
END XOR3X1H7R

MACRO XOR3X1P4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR3X1P4H7R 0 0 ;
  SIZE 4.2 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.2 1.48 ;
        RECT 3.29 1.05 3.38 1.48 ;
        RECT 2.81 1.035 2.9 1.48 ;
        RECT 1.575 1.2 1.665 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.2 0.08 ;
        RECT 3.76 -0.08 3.85 0.33 ;
        RECT 3.28 -0.08 3.37 0.345 ;
        RECT 1.59 -0.08 1.68 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.475 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.765 0.375 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.35 0.655 3.65 0.745 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.68 1.055 4.1 1.145 ;
        RECT 4.01 0.301 4.1 1.145 ;
      LAYER MET2 ;
        RECT 3.85 0.84 3.95 1.22 ;
      LAYER VIA1 ;
        RECT 3.855 1.055 3.945 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.335 0.435 2.425 1.015 ;
      RECT 3.194 0.835 3.92 0.925 ;
      RECT 3.83 0.66 3.92 0.925 ;
      RECT 3.155 0.777 3.194 0.906 ;
      RECT 3.109 0.735 3.155 0.863 ;
      RECT 3.109 0.816 3.232 0.863 ;
      RECT 3.063 0.689 3.109 0.817 ;
      RECT 3.017 0.643 3.063 0.771 ;
      RECT 2.979 0.689 3.109 0.729 ;
      RECT 2.335 0.62 3.017 0.71 ;
      RECT 2.07 0.435 2.665 0.525 ;
      RECT 2.525 0.35 2.665 0.525 ;
      RECT 2.07 0.205 2.16 0.525 ;
      RECT 2.775 0.44 3.6 0.53 ;
      RECT 3.51 0.205 3.6 0.53 ;
      RECT 2.775 0.35 2.915 0.53 ;
      RECT 2.07 1.105 2.72 1.195 ;
      RECT 2.63 0.835 2.72 1.195 ;
      RECT 3.04 0.967 3.13 1.14 ;
      RECT 2.07 1.035 2.16 1.195 ;
      RECT 3.022 0.89 3.04 1.018 ;
      RECT 2.976 0.858 3.022 0.986 ;
      RECT 2.976 0.922 3.086 0.986 ;
      RECT 2.938 0.922 3.086 0.944 ;
      RECT 2.63 0.835 2.976 0.925 ;
      RECT 3.03 0.17 3.12 0.345 ;
      RECT 2.32 0.17 2.41 0.345 ;
      RECT 2.32 0.17 3.12 0.26 ;
      RECT 1.84 0.225 1.93 1.115 ;
      RECT 1.84 0.694 2.035 0.784 ;
      RECT 0.78 1.11 1.446 1.2 ;
      RECT 0.78 1.11 1.492 1.177 ;
      RECT 1.408 1.091 1.538 1.131 ;
      RECT 0.78 0.35 0.87 1.2 ;
      RECT 1.446 1.049 1.538 1.131 ;
      RECT 1.492 1.003 1.584 1.085 ;
      RECT 1.492 1.003 1.63 1.039 ;
      RECT 1.538 0.957 1.65 1.006 ;
      RECT 1.584 0.911 1.696 0.973 ;
      RECT 1.63 0.878 1.65 1.006 ;
      RECT 1.65 0.765 1.74 0.928 ;
      RECT 0.78 0.35 0.925 0.44 ;
      RECT 1.275 0.712 1.365 1.018 ;
      RECT 1.241 0.672 1.331 0.75 ;
      RECT 1.195 0.437 1.285 0.71 ;
      RECT 1.195 0.437 1.331 0.475 ;
      RECT 1.241 0.397 1.34 0.448 ;
      RECT 1.275 0.375 1.386 0.42 ;
      RECT 1.331 0.319 1.34 0.448 ;
      RECT 1.34 0.205 1.43 0.375 ;
      RECT 1.285 0.347 1.43 0.375 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 1.015 0.84 1.16 0.93 ;
      RECT 1.015 0.17 1.105 0.93 ;
      RECT 0.045 0.445 0.64 0.535 ;
      RECT 0.55 0.17 0.64 0.535 ;
      RECT 1.015 0.17 1.18 0.345 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.55 0.17 1.18 0.26 ;
  END
END XOR3X1P4H7R

MACRO XOR3X2H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR3X2H7R 0 0 ;
  SIZE 4.4 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.4 1.48 ;
        RECT 3.96 1.24 4.1 1.48 ;
        RECT 3.29 1.05 3.38 1.48 ;
        RECT 2.81 1.035 2.9 1.48 ;
        RECT 1.575 1.2 1.665 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.4 0.08 ;
        RECT 4.24 -0.08 4.33 0.345 ;
        RECT 3.74 -0.08 3.83 0.33 ;
        RECT 3.26 -0.08 3.35 0.345 ;
        RECT 1.57 -0.08 1.66 0.33 ;
        RECT 0.32 -0.08 0.41 0.33 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.475 1.545 0.775 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.225 0.765 0.375 0.945 ;
      LAYER MET2 ;
        RECT 0.25 0.625 0.35 1.16 ;
      LAYER VIA1 ;
        RECT 0.255 0.855 0.345 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.35 0.625 3.575 0.745 ;
      LAYER MET2 ;
        RECT 3.45 0.425 3.55 0.96 ;
      LAYER VIA1 ;
        RECT 3.455 0.655 3.545 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.68 1.055 4.08 1.145 ;
        RECT 3.99 0.205 4.08 1.145 ;
      LAYER MET2 ;
        RECT 3.85 0.84 3.95 1.22 ;
      LAYER VIA1 ;
        RECT 3.855 1.055 3.945 1.145 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.335 0.435 2.425 1.015 ;
      RECT 3.194 0.835 3.895 0.925 ;
      RECT 3.805 0.785 3.895 0.925 ;
      RECT 3.155 0.777 3.194 0.906 ;
      RECT 3.109 0.735 3.155 0.863 ;
      RECT 3.109 0.816 3.232 0.863 ;
      RECT 3.063 0.689 3.109 0.817 ;
      RECT 3.017 0.643 3.063 0.771 ;
      RECT 2.979 0.689 3.109 0.729 ;
      RECT 2.335 0.62 3.017 0.71 ;
      RECT 2.05 0.435 2.645 0.525 ;
      RECT 2.505 0.35 2.645 0.525 ;
      RECT 2.05 0.205 2.14 0.525 ;
      RECT 2.755 0.44 3.58 0.53 ;
      RECT 3.49 0.205 3.58 0.53 ;
      RECT 2.755 0.35 2.895 0.53 ;
      RECT 2.07 1.14 2.72 1.23 ;
      RECT 2.63 0.835 2.72 1.23 ;
      RECT 2.07 1.035 2.16 1.23 ;
      RECT 3.04 0.967 3.13 1.135 ;
      RECT 3.022 0.89 3.04 1.018 ;
      RECT 2.976 0.858 3.022 0.986 ;
      RECT 2.976 0.922 3.086 0.986 ;
      RECT 2.938 0.922 3.086 0.944 ;
      RECT 2.63 0.835 2.976 0.925 ;
      RECT 3.01 0.17 3.1 0.345 ;
      RECT 2.3 0.17 2.39 0.345 ;
      RECT 2.3 0.17 3.1 0.26 ;
      RECT 1.84 0.255 1.93 1.075 ;
      RECT 1.84 0.694 2.035 0.784 ;
      RECT 1.82 0.255 1.93 0.395 ;
      RECT 0.78 1.14 1.416 1.23 ;
      RECT 0.78 1.14 1.462 1.207 ;
      RECT 1.378 1.121 1.508 1.161 ;
      RECT 0.78 0.35 0.87 1.23 ;
      RECT 1.416 1.079 1.508 1.161 ;
      RECT 1.462 1.033 1.554 1.115 ;
      RECT 1.508 0.987 1.6 1.069 ;
      RECT 1.508 0.987 1.646 1.023 ;
      RECT 1.554 0.941 1.66 0.993 ;
      RECT 1.6 0.895 1.706 0.963 ;
      RECT 1.646 0.865 1.66 0.993 ;
      RECT 1.66 0.725 1.75 0.918 ;
      RECT 0.78 0.35 0.925 0.44 ;
      RECT 1.275 0.712 1.365 1.018 ;
      RECT 1.241 0.396 1.285 0.75 ;
      RECT 1.241 0.672 1.331 0.75 ;
      RECT 1.195 0.436 1.285 0.71 ;
      RECT 1.285 0.351 1.32 0.48 ;
      RECT 1.275 0.374 1.366 0.439 ;
      RECT 1.32 0.205 1.41 0.394 ;
      RECT 0.045 1.04 0.185 1.13 ;
      RECT 0.045 0.23 0.135 1.13 ;
      RECT 1.015 0.84 1.16 0.93 ;
      RECT 1.015 0.17 1.105 0.93 ;
      RECT 0.045 0.445 0.64 0.535 ;
      RECT 0.55 0.17 0.64 0.535 ;
      RECT 1.015 0.17 1.18 0.345 ;
      RECT 0.045 0.23 0.185 0.32 ;
      RECT 0.55 0.17 1.18 0.26 ;
  END
END XOR3X2H7R

MACRO XOR3X3H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR3X3H7R 0 0 ;
  SIZE 4.6 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 4.6 1.48 ;
        RECT 4.435 1.035 4.525 1.48 ;
        RECT 3.863 1.195 4.003 1.48 ;
        RECT 3.338 1.195 3.478 1.48 ;
        RECT 1.603 1.2 1.693 1.48 ;
        RECT 0.32 1.07 0.41 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 4.6 0.08 ;
        RECT 4.403 -0.08 4.493 0.345 ;
        RECT 3.903 -0.08 3.993 0.345 ;
        RECT 3.313 -0.08 3.403 0.33 ;
        RECT 1.618 -0.08 1.708 0.33 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.455 0.56 1.555 0.83 ;
      LAYER MET2 ;
        RECT 1.45 0.43 1.55 0.96 ;
      LAYER VIA1 ;
        RECT 1.455 0.655 1.545 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.505 0.645 3.775 0.745 ;
      LAYER MET2 ;
        RECT 3.65 0.43 3.75 0.96 ;
      LAYER VIA1 ;
        RECT 3.655 0.655 3.745 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.143 1.06 4.345 1.15 ;
        RECT 4.255 0.471 4.345 1.15 ;
        RECT 4.199 0.426 4.301 0.497 ;
        RECT 4.153 0.397 4.255 0.452 ;
        RECT 4.243 0.471 4.345 0.525 ;
        RECT 4.153 0.285 4.243 0.452 ;
      LAYER MET2 ;
        RECT 4.25 0.425 4.35 0.96 ;
      LAYER VIA1 ;
        RECT 4.255 0.655 4.345 0.745 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.148 1.105 3.223 1.195 ;
      RECT 3.133 0.73 3.223 1.195 ;
      RECT 3.133 1.015 3.969 1.105 ;
      RECT 2.148 0.35 2.253 1.195 ;
      RECT 3.133 1.015 4.015 1.082 ;
      RECT 3.931 0.996 4.061 1.036 ;
      RECT 3.969 0.954 4.073 1.007 ;
      RECT 4.073 0.5 4.119 0.978 ;
      RECT 4.015 0.908 4.119 0.978 ;
      RECT 4.061 0.879 4.073 1.007 ;
      RECT 4.073 0.545 4.163 0.933 ;
      RECT 4.031 0.456 4.073 0.584 ;
      RECT 3.993 0.5 4.119 0.544 ;
      RECT 3.643 0.435 4.031 0.525 ;
      RECT 3.643 0.265 3.733 0.525 ;
      RECT 2.428 0.925 3.043 1.015 ;
      RECT 2.953 0.55 3.043 1.015 ;
      RECT 3.313 0.835 3.893 0.925 ;
      RECT 2.428 0.35 2.518 1.015 ;
      RECT 3.313 0.835 3.939 0.902 ;
      RECT 3.893 0.645 3.983 0.857 ;
      RECT 3.855 0.816 3.983 0.857 ;
      RECT 3.313 0.55 3.403 0.925 ;
      RECT 2.953 0.55 3.403 0.64 ;
      RECT 1.843 0.94 2.058 1.03 ;
      RECT 1.968 0.17 2.058 1.03 ;
      RECT 2.773 0.17 2.863 0.83 ;
      RECT 1.843 0.29 2.058 0.38 ;
      RECT 1.968 0.17 2.863 0.26 ;
      RECT 0.78 1.11 1.446 1.2 ;
      RECT 0.78 1.11 1.492 1.177 ;
      RECT 1.408 1.091 1.538 1.131 ;
      RECT 0.78 0.35 0.87 1.2 ;
      RECT 1.446 1.049 1.538 1.131 ;
      RECT 1.492 1.003 1.584 1.085 ;
      RECT 1.538 0.957 1.63 1.039 ;
      RECT 1.584 0.911 1.676 0.993 ;
      RECT 1.63 0.865 1.756 0.913 ;
      RECT 1.676 0.825 1.71 0.953 ;
      RECT 1.71 0.705 1.8 0.868 ;
      RECT 0.78 0.35 0.93 0.44 ;
      RECT 1.275 0.737 1.365 1.018 ;
      RECT 1.264 0.737 1.365 0.776 ;
      RECT 1.218 0.495 1.308 0.747 ;
      RECT 1.218 0.709 1.354 0.747 ;
      RECT 1.218 0.495 1.354 0.533 ;
      RECT 1.264 0.466 1.368 0.503 ;
      RECT 1.275 0.444 1.414 0.473 ;
      RECT 1.354 0.375 1.368 0.503 ;
      RECT 1.308 0.405 1.414 0.473 ;
      RECT 1.368 0.265 1.458 0.428 ;
      RECT 0.07 0.89 0.16 1.075 ;
      RECT 0.07 0.89 0.51 0.98 ;
      RECT 0.42 0.395 0.51 0.98 ;
      RECT 1.02 0.82 1.16 0.91 ;
      RECT 1.02 0.17 1.11 0.91 ;
      RECT 0.07 0.395 0.64 0.485 ;
      RECT 0.55 0.17 0.64 0.485 ;
      RECT 0.07 0.265 0.16 0.485 ;
      RECT 1.02 0.17 1.228 0.345 ;
      RECT 0.55 0.17 1.228 0.26 ;
  END
END XOR3X3H7R

MACRO XOR3X4H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR3X4H7R 0 0 ;
  SIZE 5 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5 1.48 ;
        RECT 4.782 1.035 4.872 1.48 ;
        RECT 4.282 1.035 4.372 1.48 ;
        RECT 3.482 1.24 3.622 1.48 ;
        RECT 1.832 1.2 1.922 1.48 ;
        RECT 0.295 1.08 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5 0.08 ;
        RECT 4.547 -0.08 4.637 0.33 ;
        RECT 4.047 -0.08 4.137 0.345 ;
        RECT 3.457 -0.08 3.547 0.33 ;
        RECT 1.755 -0.08 1.845 0.33 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.625 0.565 1.775 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.655 0.625 3.835 0.775 ;
      LAYER MET2 ;
        RECT 3.65 0.43 3.75 0.96 ;
      LAYER VIA1 ;
        RECT 3.655 0.655 3.745 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.438 0.455 4.887 0.545 ;
        RECT 4.797 0.255 4.887 0.545 ;
        RECT 4.532 0.455 4.622 0.93 ;
        RECT 4.343 0.436 4.476 0.472 ;
        RECT 4.343 0.414 4.438 0.472 ;
        RECT 4.433 0.455 4.887 0.543 ;
        RECT 4.297 0.389 4.433 0.427 ;
        RECT 4.387 0.455 4.887 0.517 ;
        RECT 4.297 0.26 4.387 0.427 ;
      LAYER MET2 ;
        RECT 4.65 0.225 4.75 0.76 ;
      LAYER VIA1 ;
        RECT 4.655 0.455 4.745 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.488 1.065 3.367 1.155 ;
      RECT 3.277 0.665 3.367 1.155 ;
      RECT 2.488 1.065 4.023 1.135 ;
      RECT 2.488 1.065 4.069 1.112 ;
      RECT 3.277 1.045 4.115 1.066 ;
      RECT 2.488 0.923 2.578 1.155 ;
      RECT 3.985 1.026 4.115 1.066 ;
      RECT 4.023 0.984 4.115 1.066 ;
      RECT 4.069 0.938 4.161 1.02 ;
      RECT 2.482 0.852 2.488 0.98 ;
      RECT 4.069 0.938 4.207 0.974 ;
      RECT 4.115 0.892 4.217 0.946 ;
      RECT 2.438 0.878 2.534 0.955 ;
      RECT 4.217 0.475 4.263 0.918 ;
      RECT 2.392 0.35 2.482 0.91 ;
      RECT 4.161 0.846 4.263 0.918 ;
      RECT 4.207 0.818 4.217 0.946 ;
      RECT 4.217 0.52 4.307 0.873 ;
      RECT 4.205 0.446 4.217 0.574 ;
      RECT 4.167 0.52 4.307 0.549 ;
      RECT 3.787 0.44 4.205 0.53 ;
      RECT 2.292 0.35 2.482 0.49 ;
      RECT 3.787 0.305 3.877 0.53 ;
      RECT 2.757 0.885 3.187 0.975 ;
      RECT 3.097 0.485 3.187 0.975 ;
      RECT 2.754 0.845 2.757 0.974 ;
      RECT 3.457 0.865 3.947 0.955 ;
      RECT 2.708 0.821 2.754 0.949 ;
      RECT 3.457 0.865 3.993 0.932 ;
      RECT 2.662 0.775 2.708 0.903 ;
      RECT 2.662 0.866 2.795 0.903 ;
      RECT 3.909 0.846 4.037 0.887 ;
      RECT 3.457 0.485 3.547 0.955 ;
      RECT 2.618 0.35 2.662 0.858 ;
      RECT 3.947 0.804 4.037 0.887 ;
      RECT 2.572 0.35 2.662 0.813 ;
      RECT 3.993 0.759 4.083 0.842 ;
      RECT 4.037 0.62 4.127 0.797 ;
      RECT 3.097 0.485 3.547 0.575 ;
      RECT 2.112 0.17 2.202 1.015 ;
      RECT 2.917 0.17 3.007 0.795 ;
      RECT 2.112 0.655 2.267 0.795 ;
      RECT 1.98 0.23 2.202 0.32 ;
      RECT 2.112 0.17 3.007 0.26 ;
      RECT 0.78 1.11 1.704 1.2 ;
      RECT 0.78 1.11 1.75 1.177 ;
      RECT 1.666 1.091 1.796 1.131 ;
      RECT 1.31 1.055 1.4 1.2 ;
      RECT 0.78 0.35 0.87 1.2 ;
      RECT 1.704 1.049 1.796 1.131 ;
      RECT 1.75 1.003 1.842 1.085 ;
      RECT 1.796 0.957 1.888 1.039 ;
      RECT 1.842 0.911 1.93 0.995 ;
      RECT 1.888 0.867 1.976 0.951 ;
      RECT 1.93 0.665 2.02 0.906 ;
      RECT 0.78 0.35 0.93 0.44 ;
      RECT 1.54 0.878 1.63 1.018 ;
      RECT 1.537 0.844 1.54 0.973 ;
      RECT 1.491 0.82 1.537 0.948 ;
      RECT 1.445 0.774 1.491 0.902 ;
      RECT 1.445 0.862 1.572 0.902 ;
      RECT 1.401 0.48 1.445 0.857 ;
      RECT 1.355 0.525 1.445 0.812 ;
      RECT 1.355 0.525 1.491 0.563 ;
      RECT 1.401 0.48 1.505 0.533 ;
      RECT 1.445 0.435 1.551 0.503 ;
      RECT 1.491 0.405 1.505 0.533 ;
      RECT 1.505 0.29 1.595 0.458 ;
      RECT 0.07 0.89 0.16 1.035 ;
      RECT 1.045 0.17 1.135 1.005 ;
      RECT 0.07 0.89 0.51 0.98 ;
      RECT 0.42 0.395 0.51 0.98 ;
      RECT 0.07 0.395 0.64 0.485 ;
      RECT 0.55 0.17 0.64 0.485 ;
      RECT 0.07 0.305 0.16 0.485 ;
      RECT 1.045 0.23 1.39 0.32 ;
      RECT 0.55 0.17 1.135 0.26 ;
  END
END XOR3X4H7R

MACRO XOR3X6H7R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR3X6H7R 0 0 ;
  SIZE 5 BY 1.4 ;
  SYMMETRY X Y ;
  SITE core7 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 1.32 5 1.48 ;
        RECT 4.552 0.85 4.642 1.48 ;
        RECT 3.982 1.24 4.122 1.48 ;
        RECT 3.457 1.24 3.597 1.48 ;
        RECT 1.832 1.2 1.922 1.48 ;
        RECT 0.295 1.08 0.435 1.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.08 5 0.08 ;
        RECT 4.84 -0.08 4.93 0.345 ;
        RECT 4.34 -0.08 4.43 0.33 ;
        RECT 3.812 -0.08 3.952 0.32 ;
        RECT 3.247 -0.08 3.337 0.33 ;
        RECT 1.755 -0.08 1.845 0.33 ;
        RECT 0.295 -0.08 0.435 0.305 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.625 0.565 1.775 0.745 ;
      LAYER MET2 ;
        RECT 1.65 0.43 1.75 0.96 ;
      LAYER VIA1 ;
        RECT 1.655 0.655 1.745 0.745 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.055 0.625 0.235 0.775 ;
      LAYER MET2 ;
        RECT 0.05 0.43 0.15 0.96 ;
      LAYER VIA1 ;
        RECT 0.055 0.655 0.145 0.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.637 0.61 3.787 0.79 ;
      LAYER MET2 ;
        RECT 3.65 0.43 3.75 0.96 ;
      LAYER VIA1 ;
        RECT 3.655 0.655 3.745 0.745 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.817 0.455 4.907 1.145 ;
        RECT 4.287 0.455 4.907 0.545 ;
        RECT 4.59 0.295 4.68 0.545 ;
        RECT 4.287 0.455 4.377 1.13 ;
        RECT 4.223 0.431 4.333 0.494 ;
        RECT 4.177 0.407 4.287 0.448 ;
        RECT 4.286 0.455 4.907 0.534 ;
        RECT 4.177 0.397 4.286 0.448 ;
        RECT 4.269 0.455 4.907 0.526 ;
        RECT 4.133 0.366 4.269 0.403 ;
        RECT 4.133 0.32 4.223 0.403 ;
        RECT 4.087 0.19 4.177 0.358 ;
      LAYER MET2 ;
        RECT 4.45 0.225 4.55 0.76 ;
      LAYER VIA1 ;
        RECT 4.455 0.455 4.545 0.545 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.488 1.065 3.367 1.155 ;
      RECT 3.277 0.665 3.367 1.155 ;
      RECT 4.077 0.522 4.167 1.15 ;
      RECT 3.277 1.06 4.167 1.15 ;
      RECT 2.488 0.938 2.578 1.155 ;
      RECT 2.482 0.867 2.488 0.995 ;
      RECT 2.438 0.893 2.534 0.97 ;
      RECT 2.392 0.35 2.482 0.925 ;
      RECT 4.053 0.442 4.077 0.57 ;
      RECT 4.015 0.477 4.123 0.539 ;
      RECT 3.607 0.43 4.053 0.52 ;
      RECT 2.292 0.35 2.482 0.49 ;
      RECT 3.607 0.305 3.697 0.52 ;
      RECT 2.757 0.885 3.187 0.975 ;
      RECT 3.097 0.485 3.187 0.975 ;
      RECT 2.754 0.845 2.757 0.974 ;
      RECT 3.457 0.88 3.987 0.97 ;
      RECT 3.897 0.62 3.987 0.97 ;
      RECT 2.708 0.821 2.754 0.949 ;
      RECT 2.662 0.775 2.708 0.903 ;
      RECT 2.662 0.866 2.795 0.903 ;
      RECT 3.457 0.566 3.547 0.97 ;
      RECT 2.618 0.35 2.662 0.858 ;
      RECT 2.572 0.35 2.662 0.813 ;
      RECT 3.444 0.491 3.457 0.62 ;
      RECT 3.406 0.566 3.547 0.594 ;
      RECT 3.097 0.485 3.444 0.575 ;
      RECT 3.097 0.521 3.503 0.575 ;
      RECT 2.112 0.17 2.202 1.015 ;
      RECT 2.917 0.17 3.007 0.795 ;
      RECT 2.112 0.655 2.267 0.795 ;
      RECT 1.98 0.23 2.202 0.32 ;
      RECT 2.112 0.17 3.007 0.26 ;
      RECT 0.78 1.105 1.709 1.195 ;
      RECT 0.78 1.105 1.755 1.172 ;
      RECT 1.671 1.086 1.801 1.126 ;
      RECT 1.31 1.05 1.4 1.195 ;
      RECT 0.78 0.35 0.87 1.195 ;
      RECT 1.709 1.044 1.801 1.126 ;
      RECT 1.755 0.998 1.847 1.08 ;
      RECT 1.801 0.952 1.893 1.034 ;
      RECT 1.847 0.906 1.93 0.993 ;
      RECT 1.847 0.906 1.976 0.951 ;
      RECT 1.93 0.665 2.02 0.906 ;
      RECT 1.893 0.864 2.02 0.906 ;
      RECT 0.78 0.35 0.93 0.44 ;
      RECT 1.54 0.875 1.63 1.015 ;
      RECT 1.537 0.794 1.54 0.923 ;
      RECT 1.491 0.77 1.537 0.898 ;
      RECT 1.491 0.858 1.619 0.898 ;
      RECT 1.491 0.819 1.586 0.898 ;
      RECT 1.445 0.724 1.491 0.852 ;
      RECT 1.401 0.495 1.445 0.807 ;
      RECT 1.355 0.54 1.445 0.762 ;
      RECT 1.355 0.54 1.491 0.578 ;
      RECT 1.401 0.495 1.505 0.548 ;
      RECT 1.445 0.45 1.551 0.518 ;
      RECT 1.491 0.42 1.505 0.548 ;
      RECT 1.505 0.305 1.595 0.473 ;
      RECT 0.07 0.89 0.16 1.035 ;
      RECT 1.045 0.17 1.135 1.005 ;
      RECT 0.07 0.89 0.51 0.98 ;
      RECT 0.42 0.395 0.51 0.98 ;
      RECT 0.07 0.395 0.64 0.485 ;
      RECT 0.55 0.17 0.64 0.485 ;
      RECT 0.07 0.305 0.16 0.485 ;
      RECT 1.045 0.23 1.39 0.32 ;
      RECT 0.55 0.17 1.135 0.26 ;
  END
END XOR3X6H7R

END LIBRARY
