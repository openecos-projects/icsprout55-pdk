# Copyright 2025 ICsprout Integrated Circuit Co., Ltd.
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
  LAYER LEF58_ENCLOSURE STRING ;
  LAYER LEF58_WIDTH STRING ;
  LAYER LEF58_SPACING STRING ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.001 ;
LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

LAYER ACT
  TYPE MASTERSLICE ;
END ACT

LAYER NP
  TYPE MASTERSLICE ;
END NP

LAYER PP
  TYPE MASTERSLICE ;
END PP

LAYER NW1
  TYPE MASTERSLICE ;
END NW1

LAYER POLY
  TYPE MASTERSLICE ;
END POLY

LAYER CT
  TYPE CUT ;
  SPACING 0.11 ;
  WIDTH 0.09 ;
  ENCLOSURE ABOVE 0.04 0 ;
  DCCURRENTDENSITY AVERAGE 0.29 ;
END CT

LAYER MET1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.09 ;
  OFFSET 0.1 0.1 ;
  AREA 0.042 ;
  SPACING 0.09 ;
  MAXWIDTH 10 ;
  MINENCLOSEDAREA 0.18 ;
  CAPACITANCE CPERSQDIST 0.0007630 ;
  EDGECAPACITANCE 0.0000339 ;
  RESISTANCE RPERSQ 0.1122 ;
  DCCURRENTDENSITY AVERAGE 1.5 ;
END MET1

LAYER VIA1
  TYPE CUT ;
  SPACING 0.11 ;
  WIDTH 0.09 ;
  DCCURRENTDENSITY AVERAGE 0.135 ;
END VIA1

LAYER MET2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 0.1 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  MAXWIDTH 10 ;
  MINENCLOSEDAREA 0.18 ;
  CAPACITANCE CPERSQDIST 0.0011069 ;
  EDGECAPACITANCE 0.0000391 ;
  RESISTANCE RPERSQ 0.0914 ;
  DCCURRENTDENSITY AVERAGE 1.7 ;
END MET2

LAYER VIA2
  TYPE CUT ;
  SPACING 0.11 ;
  WIDTH 0.09 ;
  DCCURRENTDENSITY AVERAGE 0.135 ;
END VIA2

LAYER MET3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 0.1 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  MAXWIDTH 10 ;
  MINENCLOSEDAREA 0.18 ;
  CAPACITANCE CPERSQDIST 0.0011069 ;
  EDGECAPACITANCE 0.0000409 ;
  RESISTANCE RPERSQ 0.0914 ;
  DCCURRENTDENSITY AVERAGE 1.7 ;
END MET3

LAYER VIA3
  TYPE CUT ;
  SPACING 0.11 ;
  WIDTH 0.09 ;
  DCCURRENTDENSITY AVERAGE 0.135 ;
END VIA3

LAYER MET4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 0.1 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  MAXWIDTH 10 ;
  MINENCLOSEDAREA 0.18 ;
  CAPACITANCE CPERSQDIST 0.0011069 ;
  EDGECAPACITANCE 0.0000409 ;
  RESISTANCE RPERSQ 0.0914 ;
  DCCURRENTDENSITY AVERAGE 1.7 ;
END MET4

LAYER VIA4
  TYPE CUT ;
  SPACING 0.11 ;
  WIDTH 0.09 ;
  ENCLOSURE BELOW 0.02 0.005 ;
  DCCURRENTDENSITY AVERAGE 0.135 ;
END VIA4

LAYER MET5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 0.1 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  MAXWIDTH 10 ;
  MINENCLOSEDAREA 0.18 ;
  CAPACITANCE CPERSQDIST 0.0006259 ;
  EDGECAPACITANCE 0.0000344 ;
  RESISTANCE RPERSQ 0.0914 ;
  DCCURRENTDENSITY AVERAGE 1.7 ;
END MET5


LAYER T4V2
  TYPE CUT ;
  SPACING 0.34 ;
  WIDTH 0.36 ;
  ENCLOSURE BELOW 0.02 0.02 ;
  DCCURRENTDENSITY AVERAGE 3.2 ;
END T4V2

LAYER T4M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.8 0.8 ;
  WIDTH 0.4 ;
  OFFSET 0.1 0.1 ;
  AREA 0.4 ;
  SPACING 0.4 ;
  MAXWIDTH 20 ;
  MINENCLOSEDAREA 0.6 ;
  CAPACITANCE CPERSQDIST 0.0001299 ;
  EDGECAPACITANCE 0.0000368 ;
  RESISTANCE RPERSQ 0.0239 ;
  DCCURRENTDENSITY AVERAGE 8.1 ;
END T4M2


LAYER RV
  TYPE CUT ;
  SPACING 3 ;
  WIDTH 3 ;
  ENCLOSURE BELOW 1.5 1.5 ;
  ENCLOSURE ABOVE 1.5 1.5 ;
END RV

LAYER RDL
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 5 5 ;
  WIDTH 3 ;
  OFFSET 0.1 0.1 ;
  SPACING 2 ;
  CAPACITANCE CPERSQDIST 0.0000574 ;
  EDGECAPACITANCE 0.0000281 ;
  RESISTANCE RPERSQ 0.0151 ;
END RDL
VIA MET2_MET1_VIA1_0 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET1 ;
		RECT -0.050 -0.085 0.050 0.085 ;
	LAYER VIA1 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET2 ;
		RECT -0.050 -0.085 0.050 0.085 ;
END MET2_MET1_VIA1_0

VIA MET2_MET1_VIA1_1 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET1 ;
		RECT -0.075 -0.075 0.075 0.075 ;
	LAYER VIA1 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET2 ;
		RECT -0.050 -0.085 0.050 0.085 ;
END MET2_MET1_VIA1_1

VIA MET2_MET1_VIA1_2 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET1 ;
		RECT -0.085 -0.050 0.085 0.050 ;
	LAYER VIA1 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET2 ;
		RECT -0.050 -0.085 0.050 0.085 ;
END MET2_MET1_VIA1_2

VIA MET2_MET1_VIA1_3 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET1 ;
		RECT -0.050 -0.085 0.050 0.085 ;
	LAYER VIA1 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET2 ;
		RECT -0.075 -0.075 0.075 0.075 ;
END MET2_MET1_VIA1_3

VIA MET2_MET1_VIA1_4 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET1 ;
		RECT -0.075 -0.075 0.075 0.075 ;
	LAYER VIA1 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET2 ;
		RECT -0.075 -0.075 0.075 0.075 ;
END MET2_MET1_VIA1_4

VIA MET2_MET1_VIA1_5 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET1 ;
		RECT -0.085 -0.050 0.085 0.050 ;
	LAYER VIA1 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET2 ;
		RECT -0.075 -0.075 0.075 0.075 ;
END MET2_MET1_VIA1_5

VIA MET2_MET1_VIA1_6 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET1 ;
		RECT -0.050 -0.085 0.050 0.085 ;
	LAYER VIA1 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET2 ;
		RECT -0.085 -0.050 0.085 0.050 ;
END MET2_MET1_VIA1_6

VIA MET2_MET1_VIA1_7 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET1 ;
		RECT -0.075 -0.075 0.075 0.075 ;
	LAYER VIA1 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET2 ;
		RECT -0.085 -0.050 0.085 0.050 ;
END MET2_MET1_VIA1_7

VIA MET2_MET1_VIA1_8 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET1 ;
		RECT -0.085 -0.050 0.085 0.050 ;
	LAYER VIA1 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET2 ;
		RECT -0.085 -0.050 0.085 0.050 ;
END MET2_MET1_VIA1_8

VIA MET3_MET2_VIA2_0 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET2 ;
		RECT -0.050 -0.085 0.050 0.085 ;
	LAYER VIA2 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET3 ;
		RECT -0.050 -0.085 0.050 0.085 ;
END MET3_MET2_VIA2_0

VIA MET3_MET2_VIA2_1 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET2 ;
		RECT -0.075 -0.075 0.075 0.075 ;
	LAYER VIA2 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET3 ;
		RECT -0.050 -0.085 0.050 0.085 ;
END MET3_MET2_VIA2_1

VIA MET3_MET2_VIA2_2 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET2 ;
		RECT -0.085 -0.050 0.085 0.050 ;
	LAYER VIA2 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET3 ;
		RECT -0.050 -0.085 0.050 0.085 ;
END MET3_MET2_VIA2_2

VIA MET3_MET2_VIA2_3 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET2 ;
		RECT -0.050 -0.085 0.050 0.085 ;
	LAYER VIA2 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET3 ;
		RECT -0.075 -0.075 0.075 0.075 ;
END MET3_MET2_VIA2_3

VIA MET3_MET2_VIA2_4 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET2 ;
		RECT -0.075 -0.075 0.075 0.075 ;
	LAYER VIA2 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET3 ;
		RECT -0.075 -0.075 0.075 0.075 ;
END MET3_MET2_VIA2_4

VIA MET3_MET2_VIA2_5 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET2 ;
		RECT -0.085 -0.050 0.085 0.050 ;
	LAYER VIA2 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET3 ;
		RECT -0.075 -0.075 0.075 0.075 ;
END MET3_MET2_VIA2_5

VIA MET3_MET2_VIA2_6 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET2 ;
		RECT -0.050 -0.085 0.050 0.085 ;
	LAYER VIA2 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET3 ;
		RECT -0.085 -0.050 0.085 0.050 ;
END MET3_MET2_VIA2_6

VIA MET3_MET2_VIA2_7 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET2 ;
		RECT -0.075 -0.075 0.075 0.075 ;
	LAYER VIA2 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET3 ;
		RECT -0.085 -0.050 0.085 0.050 ;
END MET3_MET2_VIA2_7

VIA MET3_MET2_VIA2_8 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET2 ;
		RECT -0.085 -0.050 0.085 0.050 ;
	LAYER VIA2 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET3 ;
		RECT -0.085 -0.050 0.085 0.050 ;
END MET3_MET2_VIA2_8

VIA MET4_MET3_VIA3_0 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET3 ;
		RECT -0.050 -0.085 0.050 0.085 ;
	LAYER VIA3 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET4 ;
		RECT -0.050 -0.085 0.050 0.085 ;
END MET4_MET3_VIA3_0

VIA MET4_MET3_VIA3_1 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET3 ;
		RECT -0.075 -0.075 0.075 0.075 ;
	LAYER VIA3 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET4 ;
		RECT -0.050 -0.085 0.050 0.085 ;
END MET4_MET3_VIA3_1

VIA MET4_MET3_VIA3_2 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET3 ;
		RECT -0.085 -0.050 0.085 0.050 ;
	LAYER VIA3 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET4 ;
		RECT -0.050 -0.085 0.050 0.085 ;
END MET4_MET3_VIA3_2

VIA MET4_MET3_VIA3_3 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET3 ;
		RECT -0.050 -0.085 0.050 0.085 ;
	LAYER VIA3 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET4 ;
		RECT -0.075 -0.075 0.075 0.075 ;
END MET4_MET3_VIA3_3

VIA MET4_MET3_VIA3_4 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET3 ;
		RECT -0.075 -0.075 0.075 0.075 ;
	LAYER VIA3 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET4 ;
		RECT -0.075 -0.075 0.075 0.075 ;
END MET4_MET3_VIA3_4

VIA MET4_MET3_VIA3_5 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET3 ;
		RECT -0.085 -0.050 0.085 0.050 ;
	LAYER VIA3 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET4 ;
		RECT -0.075 -0.075 0.075 0.075 ;
END MET4_MET3_VIA3_5

VIA MET4_MET3_VIA3_6 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET3 ;
		RECT -0.050 -0.085 0.050 0.085 ;
	LAYER VIA3 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET4 ;
		RECT -0.085 -0.050 0.085 0.050 ;
END MET4_MET3_VIA3_6

VIA MET4_MET3_VIA3_7 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET3 ;
		RECT -0.075 -0.075 0.075 0.075 ;
	LAYER VIA3 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET4 ;
		RECT -0.085 -0.050 0.085 0.050 ;
END MET4_MET3_VIA3_7

VIA MET4_MET3_VIA3_8 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET3 ;
		RECT -0.085 -0.050 0.085 0.050 ;
	LAYER VIA3 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET4 ;
		RECT -0.085 -0.050 0.085 0.050 ;
END MET4_MET3_VIA3_8

VIA MET5_MET4_VIA4_0 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET4 ;
		RECT -0.050 -0.085 0.050 0.085 ;
	LAYER VIA4 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET5 ;
		RECT -0.050 -0.085 0.050 0.085 ;
END MET5_MET4_VIA4_0

VIA MET5_MET4_VIA4_1 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET4 ;
		RECT -0.075 -0.075 0.075 0.075 ;
	LAYER VIA4 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET5 ;
		RECT -0.050 -0.085 0.050 0.085 ;
END MET5_MET4_VIA4_1

VIA MET5_MET4_VIA4_2 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET4 ;
		RECT -0.085 -0.050 0.085 0.050 ;
	LAYER VIA4 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET5 ;
		RECT -0.050 -0.085 0.050 0.085 ;
END MET5_MET4_VIA4_2

VIA MET5_MET4_VIA4_3 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET4 ;
		RECT -0.050 -0.085 0.050 0.085 ;
	LAYER VIA4 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET5 ;
		RECT -0.075 -0.075 0.075 0.075 ;
END MET5_MET4_VIA4_3

VIA MET5_MET4_VIA4_4 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET4 ;
		RECT -0.075 -0.075 0.075 0.075 ;
	LAYER VIA4 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET5 ;
		RECT -0.075 -0.075 0.075 0.075 ;
END MET5_MET4_VIA4_4

VIA MET5_MET4_VIA4_5 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET4 ;
		RECT -0.085 -0.050 0.085 0.050 ;
	LAYER VIA4 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET5 ;
		RECT -0.075 -0.075 0.075 0.075 ;
END MET5_MET4_VIA4_5

VIA MET5_MET4_VIA4_6 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET4 ;
		RECT -0.050 -0.085 0.050 0.085 ;
	LAYER VIA4 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET5 ;
		RECT -0.085 -0.050 0.085 0.050 ;
END MET5_MET4_VIA4_6

VIA MET5_MET4_VIA4_7 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET4 ;
		RECT -0.075 -0.075 0.075 0.075 ;
	LAYER VIA4 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET5 ;
		RECT -0.085 -0.050 0.085 0.050 ;
END MET5_MET4_VIA4_7

VIA MET5_MET4_VIA4_8 DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER MET4 ;
		RECT -0.085 -0.050 0.085 0.050 ;
	LAYER VIA4 ;
		RECT -0.045 -0.045 0.045 0.045 ;
	LAYER MET5 ;
		RECT -0.085 -0.050 0.085 0.050 ;
END MET5_MET4_VIA4_8


VIA T4M2_MET5 DEFAULT
    RESISTANCE 2.5000000000 ;
    LAYER MET5 ;
        RECT -0.19 -0.23  0.19  0.23 ;
    LAYER T4V2 ;
        RECT -0.18 -0.18 0.18  0.18 ;
    LAYER T4M2 ;
        RECT -0.2 -0.2  0.2  0.2 ;
END T4M2_MET5

VIA RDL_T4M2 DEFAULT
    RESISTANCE 2.5000000000 ;
    LAYER T4M2 ;
        RECT -3 -3  3  3 ;
    LAYER RV ;
        RECT -1.5 -1.5 1.5  1.5 ;
    LAYER RDL ;
        RECT -3 -3  3  3 ;
END RDL_T4M2


VIARULE MET2_MET1 GENERATE DEFAULT
  LAYER MET1 ;
    ENCLOSURE 0.04 0 ;
  LAYER MET2 ;
    ENCLOSURE 0.04 0.005 ;
  LAYER VIA1 ;
    RECT -0.045 -0.045 0.045 0.045 ;
    SPACING 0.13 BY 0.13 ;
END MET2_MET1

VIARULE MET3_MET2 GENERATE DEFAULT
  LAYER MET2 ;
    ENCLOSURE 0.04 0.005 ;
  LAYER MET3 ;
    ENCLOSURE 0.04 0.005 ;
  LAYER VIA2 ;
    RECT -0.045 -0.045 0.045 0.045 ;
    SPACING 0.13 BY 0.13 ;
END MET3_MET2

VIARULE MET4_MET3 GENERATE DEFAULT
  LAYER MET3 ;
    ENCLOSURE 0.04 0.005 ;
  LAYER MET4 ;
    ENCLOSURE 0.04 0.005 ;
  LAYER VIA3 ;
    RECT -0.045 -0.045 0.045 0.045 ;
    SPACING 0.13 BY 0.13 ;
END MET4_MET3

VIARULE MET5_MET4 GENERATE DEFAULT
  LAYER MET4 ;
    ENCLOSURE 0.04 0.005 ;
  LAYER MET5 ;
    ENCLOSURE 0.04 0.005 ;
  LAYER VIA4 ;
    RECT -0.045 -0.045 0.045 0.045 ;
    SPACING 0.13 BY 0.13 ;
END MET5_MET4

VIARULE T4M2_MET5 GENERATE DEFAULT
  LAYER MET5 ;
    ENCLOSURE 0.1 0.05 ;
  LAYER T4M2 ;
    ENCLOSURE 0.5 0.02 ;
  LAYER T4V2 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 1 BY 1 ;
END T4M2_MET5

VIARULE RDL_T4M2 GENERATE DEFAULT
  LAYER T4M2 ;
    ENCLOSURE 1.5 1.5 ;
  LAYER RV ;
    ENCLOSURE 1.5 1.5 ;
  LAYER RDL ;
    RECT -1.5 -1.5 1.5 1.5 ;
    SPACING 6 BY 6 ;
END RDL_T4M2

NONDEFAULTRULE virtuosoDefaultTaper
  LAYER POLY
    WIDTH 0.06 ;
  END POLY
  LAYER MET1
    WIDTH 0.09 ;
  END MET1
  USEVIARULE MET1_POLY ;
END virtuosoDefaultTaper

SITE CoreSite
    SIZE 0.2 BY 1.4 ;
    SYMMETRY Y ;
    CLASS CORE ;
END CoreSite

SITE core7
    SIZE 0.200 BY 1.400 ;
    CLASS CORE ;
    SYMMETRY Y  ;
END core7

SITE core9
    SIZE 0.200 BY 1.800 ;
    CLASS CORE ;
    SYMMETRY Y  ;
END core9

END LIBRARY